`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 05/12/2021 11:02:02 PM
// Design Name: 
// Module Name: mux_2i1o_256b_dly
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module mux_2i1O_256b_dly(
    input  clk_i,
    input  ce_i,

    input  sel_i,
    input  [255:0] in_0_i,
    input  [255:0] in_1_i,

    output [255:0] out_o
    );
    wire   [255:0] out;

   LUT3 #(
         .INIT(8'hca)         // Specify LUT Contents
         )mux_255(.O(out[255]),     // LUT general output
            .I0(in_0_i[255]), // LUT input
            .I1(in_1_i[255]), // LUT input
            .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_254(.O(out[254]),     // LUT general output
                    .I0(in_0_i[254]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_253(.O(out[253]),     // LUT general output
                    .I0(in_0_i[253]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_252(.O(out[252]),     // LUT general output
                    .I0(in_0_i[252]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_251(.O(out[251]),     // LUT general output
                    .I0(in_0_i[251]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_250(.O(out[250]),     // LUT general output
                    .I0(in_0_i[250]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_249(.O(out[249]),     // LUT general output
                    .I0(in_0_i[249]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_248(.O(out[248]),     // LUT general output
                    .I0(in_0_i[248]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_247(.O(out[247]),     // LUT general output
                    .I0(in_0_i[247]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_246(.O(out[246]),     // LUT general output
                    .I0(in_0_i[246]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_245(.O(out[245]),     // LUT general output
                    .I0(in_0_i[245]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_244(.O(out[244]),     // LUT general output
                    .I0(in_0_i[244]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_243(.O(out[243]),     // LUT general output
                    .I0(in_0_i[243]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_242(.O(out[242]),     // LUT general output
                    .I0(in_0_i[242]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_241(.O(out[241]),     // LUT general output
                    .I0(in_0_i[241]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_240(.O(out[240]),     // LUT general output
                    .I0(in_0_i[240]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_239(.O(out[239]),     // LUT general output
                    .I0(in_0_i[239]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_238(.O(out[238]),     // LUT general output
                    .I0(in_0_i[238]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_237(.O(out[237]),     // LUT general output
                    .I0(in_0_i[237]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_236(.O(out[236]),     // LUT general output
                    .I0(in_0_i[236]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_235(.O(out[235]),     // LUT general output
                    .I0(in_0_i[235]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_234(.O(out[234]),     // LUT general output
                    .I0(in_0_i[234]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_233(.O(out[233]),     // LUT general output
                    .I0(in_0_i[233]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_232(.O(out[232]),     // LUT general output
                    .I0(in_0_i[232]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_231(.O(out[231]),     // LUT general output
                    .I0(in_0_i[231]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_230(.O(out[230]),     // LUT general output
                    .I0(in_0_i[230]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_229(.O(out[229]),     // LUT general output
                    .I0(in_0_i[229]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_228(.O(out[228]),     // LUT general output
                    .I0(in_0_i[228]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_227(.O(out[227]),     // LUT general output
                    .I0(in_0_i[227]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_226(.O(out[226]),     // LUT general output
                    .I0(in_0_i[226]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_225(.O(out[225]),     // LUT general output
                    .I0(in_0_i[225]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_224(.O(out[224]),     // LUT general output
                    .I0(in_0_i[224]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_223(.O(out[223]),     // LUT general output
                    .I0(in_0_i[223]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_222(.O(out[222]),     // LUT general output
                    .I0(in_0_i[222]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_221(.O(out[221]),     // LUT general output
                    .I0(in_0_i[221]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_220(.O(out[220]),     // LUT general output
                    .I0(in_0_i[220]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_219(.O(out[219]),     // LUT general output
                    .I0(in_0_i[219]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_218(.O(out[218]),     // LUT general output
                    .I0(in_0_i[218]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_217(.O(out[217]),     // LUT general output
                    .I0(in_0_i[217]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_216(.O(out[216]),     // LUT general output
                    .I0(in_0_i[216]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_215(.O(out[215]),     // LUT general output
                    .I0(in_0_i[215]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_214(.O(out[214]),     // LUT general output
                    .I0(in_0_i[214]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_213(.O(out[213]),     // LUT general output
                    .I0(in_0_i[213]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_212(.O(out[212]),     // LUT general output
                    .I0(in_0_i[212]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_211(.O(out[211]),     // LUT general output
                    .I0(in_0_i[211]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_210(.O(out[210]),     // LUT general output
                    .I0(in_0_i[210]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_209(.O(out[209]),     // LUT general output
                    .I0(in_0_i[209]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_208(.O(out[208]),     // LUT general output
                    .I0(in_0_i[208]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_207(.O(out[207]),     // LUT general output
                    .I0(in_0_i[207]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_206(.O(out[206]),     // LUT general output
                    .I0(in_0_i[206]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_205(.O(out[205]),     // LUT general output
                    .I0(in_0_i[205]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_204(.O(out[204]),     // LUT general output
                    .I0(in_0_i[204]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_203(.O(out[203]),     // LUT general output
                    .I0(in_0_i[203]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_202(.O(out[202]),     // LUT general output
                    .I0(in_0_i[202]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_201(.O(out[201]),     // LUT general output
                    .I0(in_0_i[201]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_200(.O(out[200]),     // LUT general output
                    .I0(in_0_i[200]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_199(.O(out[199]),     // LUT general output
                    .I0(in_0_i[199]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_198(.O(out[198]),     // LUT general output
                    .I0(in_0_i[198]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_197(.O(out[197]),     // LUT general output
                    .I0(in_0_i[197]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_196(.O(out[196]),     // LUT general output
                    .I0(in_0_i[196]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_195(.O(out[195]),     // LUT general output
                    .I0(in_0_i[195]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_194(.O(out[194]),     // LUT general output
                    .I0(in_0_i[194]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_193(.O(out[193]),     // LUT general output
                    .I0(in_0_i[193]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_192(.O(out[192]),     // LUT general output
                    .I0(in_0_i[192]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_191(.O(out[191]),     // LUT general output
                    .I0(in_0_i[191]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_190(.O(out[190]),     // LUT general output
                    .I0(in_0_i[190]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_189(.O(out[189]),     // LUT general output
                    .I0(in_0_i[189]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_188(.O(out[188]),     // LUT general output
                    .I0(in_0_i[188]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_187(.O(out[187]),     // LUT general output
                    .I0(in_0_i[187]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_186(.O(out[186]),     // LUT general output
                    .I0(in_0_i[186]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_185(.O(out[185]),     // LUT general output
                    .I0(in_0_i[185]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_184(.O(out[184]),     // LUT general output
                    .I0(in_0_i[184]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_183(.O(out[183]),     // LUT general output
                    .I0(in_0_i[183]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_182(.O(out[182]),     // LUT general output
                    .I0(in_0_i[182]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_181(.O(out[181]),     // LUT general output
                    .I0(in_0_i[181]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_180(.O(out[180]),     // LUT general output
                    .I0(in_0_i[180]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_179(.O(out[179]),     // LUT general output
                    .I0(in_0_i[179]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_178(.O(out[178]),     // LUT general output
                    .I0(in_0_i[178]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_177(.O(out[177]),     // LUT general output
                    .I0(in_0_i[177]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_176(.O(out[176]),     // LUT general output
                    .I0(in_0_i[176]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_175(.O(out[175]),     // LUT general output
                    .I0(in_0_i[175]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_174(.O(out[174]),     // LUT general output
                    .I0(in_0_i[174]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_173(.O(out[173]),     // LUT general output
                    .I0(in_0_i[173]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_172(.O(out[172]),     // LUT general output
                    .I0(in_0_i[172]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_171(.O(out[171]),     // LUT general output
                    .I0(in_0_i[171]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_170(.O(out[170]),     // LUT general output
                    .I0(in_0_i[170]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_169(.O(out[169]),     // LUT general output
                    .I0(in_0_i[169]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_168(.O(out[168]),     // LUT general output
                    .I0(in_0_i[168]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_167(.O(out[167]),     // LUT general output
                    .I0(in_0_i[167]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_166(.O(out[166]),     // LUT general output
                    .I0(in_0_i[166]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_165(.O(out[165]),     // LUT general output
                    .I0(in_0_i[165]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_164(.O(out[164]),     // LUT general output
                    .I0(in_0_i[164]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_163(.O(out[163]),     // LUT general output
                    .I0(in_0_i[163]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_162(.O(out[162]),     // LUT general output
                    .I0(in_0_i[162]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_161(.O(out[161]),     // LUT general output
                    .I0(in_0_i[161]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_160(.O(out[160]),     // LUT general output
                    .I0(in_0_i[160]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_159(.O(out[159]),     // LUT general output
                    .I0(in_0_i[159]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_158(.O(out[158]),     // LUT general output
                    .I0(in_0_i[158]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_157(.O(out[157]),     // LUT general output
                    .I0(in_0_i[157]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_156(.O(out[156]),     // LUT general output
                    .I0(in_0_i[156]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_155(.O(out[155]),     // LUT general output
                    .I0(in_0_i[155]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_154(.O(out[154]),     // LUT general output
                    .I0(in_0_i[154]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_153(.O(out[153]),     // LUT general output
                    .I0(in_0_i[153]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_152(.O(out[152]),     // LUT general output
                    .I0(in_0_i[152]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_151(.O(out[151]),     // LUT general output
                    .I0(in_0_i[151]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_150(.O(out[150]),     // LUT general output
                    .I0(in_0_i[150]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_149(.O(out[149]),     // LUT general output
                    .I0(in_0_i[149]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_148(.O(out[148]),     // LUT general output
                    .I0(in_0_i[148]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_147(.O(out[147]),     // LUT general output
                    .I0(in_0_i[147]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_146(.O(out[146]),     // LUT general output
                    .I0(in_0_i[146]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_145(.O(out[145]),     // LUT general output
                    .I0(in_0_i[145]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_144(.O(out[144]),     // LUT general output
                    .I0(in_0_i[144]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_143(.O(out[143]),     // LUT general output
                    .I0(in_0_i[143]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_142(.O(out[142]),     // LUT general output
                    .I0(in_0_i[142]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_141(.O(out[141]),     // LUT general output
                    .I0(in_0_i[141]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_140(.O(out[140]),     // LUT general output
                    .I0(in_0_i[140]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_139(.O(out[139]),     // LUT general output
                    .I0(in_0_i[139]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_138(.O(out[138]),     // LUT general output
                    .I0(in_0_i[138]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_137(.O(out[137]),     // LUT general output
                    .I0(in_0_i[137]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_136(.O(out[136]),     // LUT general output
                    .I0(in_0_i[136]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_135(.O(out[135]),     // LUT general output
                    .I0(in_0_i[135]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_134(.O(out[134]),     // LUT general output
                    .I0(in_0_i[134]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_133(.O(out[133]),     // LUT general output
                    .I0(in_0_i[133]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_132(.O(out[132]),     // LUT general output
                    .I0(in_0_i[132]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_131(.O(out[131]),     // LUT general output
                    .I0(in_0_i[131]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_130(.O(out[130]),     // LUT general output
                    .I0(in_0_i[130]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_129(.O(out[129]),     // LUT general output
                    .I0(in_0_i[129]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_128(.O(out[128]),     // LUT general output
                    .I0(in_0_i[128]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_127(.O(out[127]),     // LUT general output
                    .I0(in_0_i[127]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_126(.O(out[126]),     // LUT general output
                    .I0(in_0_i[126]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_125(.O(out[125]),     // LUT general output
                    .I0(in_0_i[125]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_124(.O(out[124]),     // LUT general output
                    .I0(in_0_i[124]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_123(.O(out[123]),     // LUT general output
                    .I0(in_0_i[123]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_122(.O(out[122]),     // LUT general output
                    .I0(in_0_i[122]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_121(.O(out[121]),     // LUT general output
                    .I0(in_0_i[121]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_120(.O(out[120]),     // LUT general output
                    .I0(in_0_i[120]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_119(.O(out[119]),     // LUT general output
                    .I0(in_0_i[119]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_118(.O(out[118]),     // LUT general output
                    .I0(in_0_i[118]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_117(.O(out[117]),     // LUT general output
                    .I0(in_0_i[117]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_116(.O(out[116]),     // LUT general output
                    .I0(in_0_i[116]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_115(.O(out[115]),     // LUT general output
                    .I0(in_0_i[115]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_114(.O(out[114]),     // LUT general output
                    .I0(in_0_i[114]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_113(.O(out[113]),     // LUT general output
                    .I0(in_0_i[113]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_112(.O(out[112]),     // LUT general output
                    .I0(in_0_i[112]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_111(.O(out[111]),     // LUT general output
                    .I0(in_0_i[111]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_110(.O(out[110]),     // LUT general output
                    .I0(in_0_i[110]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_109(.O(out[109]),     // LUT general output
                    .I0(in_0_i[109]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_108(.O(out[108]),     // LUT general output
                    .I0(in_0_i[108]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_107(.O(out[107]),     // LUT general output
                    .I0(in_0_i[107]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_106(.O(out[106]),     // LUT general output
                    .I0(in_0_i[106]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_105(.O(out[105]),     // LUT general output
                    .I0(in_0_i[105]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_104(.O(out[104]),     // LUT general output
                    .I0(in_0_i[104]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_103(.O(out[103]),     // LUT general output
                    .I0(in_0_i[103]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_102(.O(out[102]),     // LUT general output
                    .I0(in_0_i[102]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_101(.O(out[101]),     // LUT general output
                    .I0(in_0_i[101]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_100(.O(out[100]),     // LUT general output
                    .I0(in_0_i[100]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_99(.O(out[99]),     // LUT general output
                    .I0(in_0_i[99]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_98(.O(out[98]),     // LUT general output
                    .I0(in_0_i[98]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_97(.O(out[97]),     // LUT general output
                    .I0(in_0_i[97]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_96(.O(out[96]),     // LUT general output
                    .I0(in_0_i[96]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_95(.O(out[95]),     // LUT general output
                    .I0(in_0_i[95]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_94(.O(out[94]),     // LUT general output
                    .I0(in_0_i[94]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_93(.O(out[93]),     // LUT general output
                    .I0(in_0_i[93]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_92(.O(out[92]),     // LUT general output
                    .I0(in_0_i[92]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_91(.O(out[91]),     // LUT general output
                    .I0(in_0_i[91]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_90(.O(out[90]),     // LUT general output
                    .I0(in_0_i[90]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_89(.O(out[89]),     // LUT general output
                    .I0(in_0_i[89]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_88(.O(out[88]),     // LUT general output
                    .I0(in_0_i[88]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_87(.O(out[87]),     // LUT general output
                    .I0(in_0_i[87]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_86(.O(out[86]),     // LUT general output
                    .I0(in_0_i[86]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_85(.O(out[85]),     // LUT general output
                    .I0(in_0_i[85]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_84(.O(out[84]),     // LUT general output
                    .I0(in_0_i[84]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_83(.O(out[83]),     // LUT general output
                    .I0(in_0_i[83]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_82(.O(out[82]),     // LUT general output
                    .I0(in_0_i[82]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_81(.O(out[81]),     // LUT general output
                    .I0(in_0_i[81]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_80(.O(out[80]),     // LUT general output
                    .I0(in_0_i[80]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_79(.O(out[79]),     // LUT general output
                    .I0(in_0_i[79]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_78(.O(out[78]),     // LUT general output
                    .I0(in_0_i[78]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_77(.O(out[77]),     // LUT general output
                    .I0(in_0_i[77]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_76(.O(out[76]),     // LUT general output
                    .I0(in_0_i[76]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_75(.O(out[75]),     // LUT general output
                    .I0(in_0_i[75]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_74(.O(out[74]),     // LUT general output
                    .I0(in_0_i[74]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_73(.O(out[73]),     // LUT general output
                    .I0(in_0_i[73]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_72(.O(out[72]),     // LUT general output
                    .I0(in_0_i[72]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_71(.O(out[71]),     // LUT general output
                    .I0(in_0_i[71]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_70(.O(out[70]),     // LUT general output
                    .I0(in_0_i[70]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_69(.O(out[69]),     // LUT general output
                    .I0(in_0_i[69]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_68(.O(out[68]),     // LUT general output
                    .I0(in_0_i[68]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_67(.O(out[67]),     // LUT general output
                    .I0(in_0_i[67]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_66(.O(out[66]),     // LUT general output
                    .I0(in_0_i[66]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_65(.O(out[65]),     // LUT general output
                    .I0(in_0_i[65]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_64(.O(out[64]),     // LUT general output
                    .I0(in_0_i[64]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_63(.O(out[63]),     // LUT general output
                    .I0(in_0_i[63]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_62(.O(out[62]),     // LUT general output
                    .I0(in_0_i[62]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_61(.O(out[61]),     // LUT general output
                    .I0(in_0_i[61]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_60(.O(out[60]),     // LUT general output
                    .I0(in_0_i[60]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_59(.O(out[59]),     // LUT general output
                    .I0(in_0_i[59]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_58(.O(out[58]),     // LUT general output
                    .I0(in_0_i[58]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_57(.O(out[57]),     // LUT general output
                    .I0(in_0_i[57]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_56(.O(out[56]),     // LUT general output
                    .I0(in_0_i[56]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_55(.O(out[55]),     // LUT general output
                    .I0(in_0_i[55]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_54(.O(out[54]),     // LUT general output
                    .I0(in_0_i[54]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_53(.O(out[53]),     // LUT general output
                    .I0(in_0_i[53]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_52(.O(out[52]),     // LUT general output
                    .I0(in_0_i[52]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_51(.O(out[51]),     // LUT general output
                    .I0(in_0_i[51]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_50(.O(out[50]),     // LUT general output
                    .I0(in_0_i[50]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_49(.O(out[49]),     // LUT general output
                    .I0(in_0_i[49]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_48(.O(out[48]),     // LUT general output
                    .I0(in_0_i[48]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_47(.O(out[47]),     // LUT general output
                    .I0(in_0_i[47]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_46(.O(out[46]),     // LUT general output
                    .I0(in_0_i[46]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_45(.O(out[45]),     // LUT general output
                    .I0(in_0_i[45]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_44(.O(out[44]),     // LUT general output
                    .I0(in_0_i[44]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_43(.O(out[43]),     // LUT general output
                    .I0(in_0_i[43]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_42(.O(out[42]),     // LUT general output
                    .I0(in_0_i[42]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_41(.O(out[41]),     // LUT general output
                    .I0(in_0_i[41]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_40(.O(out[40]),     // LUT general output
                    .I0(in_0_i[40]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_39(.O(out[39]),     // LUT general output
                    .I0(in_0_i[39]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_38(.O(out[38]),     // LUT general output
                    .I0(in_0_i[38]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_37(.O(out[37]),     // LUT general output
                    .I0(in_0_i[37]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_36(.O(out[36]),     // LUT general output
                    .I0(in_0_i[36]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_35(.O(out[35]),     // LUT general output
                    .I0(in_0_i[35]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_34(.O(out[34]),     // LUT general output
                    .I0(in_0_i[34]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_33(.O(out[33]),     // LUT general output
                    .I0(in_0_i[33]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_32(.O(out[32]),     // LUT general output
                    .I0(in_0_i[32]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_31(.O(out[31]),     // LUT general output
                    .I0(in_0_i[31]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_30(.O(out[30]),     // LUT general output
                    .I0(in_0_i[30]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_29(.O(out[29]),     // LUT general output
                    .I0(in_0_i[29]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_28(.O(out[28]),     // LUT general output
                    .I0(in_0_i[28]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_27(.O(out[27]),     // LUT general output
                    .I0(in_0_i[27]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_26(.O(out[26]),     // LUT general output
                    .I0(in_0_i[26]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_25(.O(out[25]),     // LUT general output
                    .I0(in_0_i[25]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_24(.O(out[24]),     // LUT general output
                    .I0(in_0_i[24]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_23(.O(out[23]),     // LUT general output
                    .I0(in_0_i[23]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_22(.O(out[22]),     // LUT general output
                    .I0(in_0_i[22]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_21(.O(out[21]),     // LUT general output
                    .I0(in_0_i[21]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_20(.O(out[20]),     // LUT general output
                    .I0(in_0_i[20]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_19(.O(out[19]),     // LUT general output
                    .I0(in_0_i[19]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_18(.O(out[18]),     // LUT general output
                    .I0(in_0_i[18]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_17(.O(out[17]),     // LUT general output
                    .I0(in_0_i[17]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_16(.O(out[16]),     // LUT general output
                    .I0(in_0_i[16]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_15(.O(out[15]),     // LUT general output
                    .I0(in_0_i[15]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_14(.O(out[14]),     // LUT general output
                    .I0(in_0_i[14]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_13(.O(out[13]),     // LUT general output
                    .I0(in_0_i[13]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_12(.O(out[12]),     // LUT general output
                    .I0(in_0_i[12]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_11(.O(out[11]),     // LUT general output
                    .I0(in_0_i[11]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_10(.O(out[10]),     // LUT general output
                    .I0(in_0_i[10]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_9(.O(out[9]),     // LUT general output
                    .I0(in_0_i[9]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_8(.O(out[8]),     // LUT general output
                    .I0(in_0_i[8]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_7(.O(out[7]),     // LUT general output
                    .I0(in_0_i[7]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_6(.O(out[6]),     // LUT general output
                    .I0(in_0_i[6]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_5(.O(out[5]),     // LUT general output
                    .I0(in_0_i[5]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_4(.O(out[4]),     // LUT general output
                    .I0(in_0_i[4]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_3(.O(out[3]),     // LUT general output
                    .I0(in_0_i[3]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_2(.O(out[2]),     // LUT general output
                    .I0(in_0_i[2]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_1(.O(out[1]),     // LUT general output
                    .I0(in_0_i[1]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );
      LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_0(.O(out[0]),     // LUT general output
                    .I0(in_0_i[0]), // LUT input
                    .I1(in_1_i[255]), // LUT input
                    .I2(sel_i)     // LUT input
          );

       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_255 (
      .Q(out_o[255]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[255])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_254 (
      .Q(out_o[254]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[254])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_253 (
      .Q(out_o[253]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[253])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_252 (
      .Q(out_o[252]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[252])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_251 (
      .Q(out_o[251]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[251])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_250 (
      .Q(out_o[250]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[250])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_249 (
      .Q(out_o[249]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[249])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_248 (
      .Q(out_o[248]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[248])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_247 (
      .Q(out_o[247]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[247])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_246 (
      .Q(out_o[246]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[246])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_245 (
      .Q(out_o[245]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[245])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_244 (
      .Q(out_o[244]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[244])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_243 (
      .Q(out_o[243]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[243])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_242 (
      .Q(out_o[242]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[242])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_241 (
      .Q(out_o[241]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[241])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_240 (
      .Q(out_o[240]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[240])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_239 (
      .Q(out_o[239]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[239])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_238 (
      .Q(out_o[238]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[238])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_237 (
      .Q(out_o[237]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[237])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_236 (
      .Q(out_o[236]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[236])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_235 (
      .Q(out_o[235]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[235])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_234 (
      .Q(out_o[234]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[234])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_233 (
      .Q(out_o[233]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[233])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_232 (
      .Q(out_o[232]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[232])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_231 (
      .Q(out_o[231]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[231])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_230 (
      .Q(out_o[230]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[230])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_229 (
      .Q(out_o[229]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[229])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_228 (
      .Q(out_o[228]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[228])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_227 (
      .Q(out_o[227]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[227])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_226 (
      .Q(out_o[226]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[226])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_225 (
      .Q(out_o[225]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[225])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_224 (
      .Q(out_o[224]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[224])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_223 (
      .Q(out_o[223]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[223])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_222 (
      .Q(out_o[222]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[222])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_221 (
      .Q(out_o[221]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[221])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_220 (
      .Q(out_o[220]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[220])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_219 (
      .Q(out_o[219]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[219])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_218 (
      .Q(out_o[218]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[218])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_217 (
      .Q(out_o[217]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[217])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_216 (
      .Q(out_o[216]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[216])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_215 (
      .Q(out_o[215]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[215])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_214 (
      .Q(out_o[214]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[214])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_213 (
      .Q(out_o[213]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[213])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_212 (
      .Q(out_o[212]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[212])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_211 (
      .Q(out_o[211]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[211])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_210 (
      .Q(out_o[210]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[210])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_209 (
      .Q(out_o[209]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[209])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_208 (
      .Q(out_o[208]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[208])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_207 (
      .Q(out_o[207]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[207])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_206 (
      .Q(out_o[206]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[206])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_205 (
      .Q(out_o[205]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[205])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_204 (
      .Q(out_o[204]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[204])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_203 (
      .Q(out_o[203]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[203])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_202 (
      .Q(out_o[202]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[202])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_201 (
      .Q(out_o[201]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[201])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_200 (
      .Q(out_o[200]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[200])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_199 (
      .Q(out_o[199]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[199])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_198 (
      .Q(out_o[198]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[198])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_197 (
      .Q(out_o[197]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[197])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_196 (
      .Q(out_o[196]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[196])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_195 (
      .Q(out_o[195]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[195])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_194 (
      .Q(out_o[194]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[194])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_193 (
      .Q(out_o[193]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[193])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_192 (
      .Q(out_o[192]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[192])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_191 (
      .Q(out_o[191]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[191])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_190 (
      .Q(out_o[190]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[190])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_189 (
      .Q(out_o[189]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[189])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_188 (
      .Q(out_o[188]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[188])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_187 (
      .Q(out_o[187]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[187])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_186 (
      .Q(out_o[186]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[186])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_185 (
      .Q(out_o[185]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[185])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_184 (
      .Q(out_o[184]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[184])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_183 (
      .Q(out_o[183]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[183])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_182 (
      .Q(out_o[182]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[182])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_181 (
      .Q(out_o[181]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[181])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_180 (
      .Q(out_o[180]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[180])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_179 (
      .Q(out_o[179]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[179])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_178 (
      .Q(out_o[178]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[178])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_177 (
      .Q(out_o[177]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[177])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_176 (
      .Q(out_o[176]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[176])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_175 (
      .Q(out_o[175]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[175])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_174 (
      .Q(out_o[174]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[174])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_173 (
      .Q(out_o[173]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[173])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_172 (
      .Q(out_o[172]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[172])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_171 (
      .Q(out_o[171]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[171])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_170 (
      .Q(out_o[170]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[170])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_169 (
      .Q(out_o[169]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[169])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_168 (
      .Q(out_o[168]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[168])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_167 (
      .Q(out_o[167]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[167])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_166 (
      .Q(out_o[166]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[166])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_165 (
      .Q(out_o[165]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[165])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_164 (
      .Q(out_o[164]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[164])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_163 (
      .Q(out_o[163]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[163])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_162 (
      .Q(out_o[162]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[162])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_161 (
      .Q(out_o[161]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[161])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_160 (
      .Q(out_o[160]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[160])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_159 (
      .Q(out_o[159]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[159])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_158 (
      .Q(out_o[158]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[158])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_157 (
      .Q(out_o[157]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[157])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_156 (
      .Q(out_o[156]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[156])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_155 (
      .Q(out_o[155]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[155])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_154 (
      .Q(out_o[154]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[154])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_153 (
      .Q(out_o[153]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[153])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_152 (
      .Q(out_o[152]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[152])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_151 (
      .Q(out_o[151]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[151])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_150 (
      .Q(out_o[150]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[150])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_149 (
      .Q(out_o[149]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[149])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_148 (
      .Q(out_o[148]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[148])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_147 (
      .Q(out_o[147]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[147])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_146 (
      .Q(out_o[146]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[146])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_145 (
      .Q(out_o[145]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[145])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_144 (
      .Q(out_o[144]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[144])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_143 (
      .Q(out_o[143]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[143])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_142 (
      .Q(out_o[142]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[142])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_141 (
      .Q(out_o[141]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[141])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_140 (
      .Q(out_o[140]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[140])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_139 (
      .Q(out_o[139]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[139])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_138 (
      .Q(out_o[138]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[138])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_137 (
      .Q(out_o[137]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[137])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_136 (
      .Q(out_o[136]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[136])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_135 (
      .Q(out_o[135]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[135])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_134 (
      .Q(out_o[134]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[134])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_133 (
      .Q(out_o[133]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[133])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_132 (
      .Q(out_o[132]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[132])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_131 (
      .Q(out_o[131]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[131])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_130 (
      .Q(out_o[130]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[130])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_129 (
      .Q(out_o[129]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[129])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_128 (
      .Q(out_o[128]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[128])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_127 (
      .Q(out_o[127]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[127])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_126 (
      .Q(out_o[126]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[126])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_125 (
      .Q(out_o[125]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[125])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_124 (
      .Q(out_o[124]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[124])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_123 (
      .Q(out_o[123]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[123])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_122 (
      .Q(out_o[122]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[122])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_121 (
      .Q(out_o[121]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[121])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_120 (
      .Q(out_o[120]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[120])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_119 (
      .Q(out_o[119]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[119])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_118 (
      .Q(out_o[118]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[118])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_117 (
      .Q(out_o[117]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[117])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_116 (
      .Q(out_o[116]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[116])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_115 (
      .Q(out_o[115]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[115])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_114 (
      .Q(out_o[114]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[114])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_113 (
      .Q(out_o[113]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[113])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_112 (
      .Q(out_o[112]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[112])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_111 (
      .Q(out_o[111]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[111])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_110 (
      .Q(out_o[110]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[110])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_109 (
      .Q(out_o[109]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[109])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_108 (
      .Q(out_o[108]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[108])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_107 (
      .Q(out_o[107]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[107])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_106 (
      .Q(out_o[106]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[106])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_105 (
      .Q(out_o[105]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[105])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_104 (
      .Q(out_o[104]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[104])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_103 (
      .Q(out_o[103]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[103])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_102 (
      .Q(out_o[102]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[102])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_101 (
      .Q(out_o[101]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[101])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_100 (
      .Q(out_o[100]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[100])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_99 (
      .Q(out_o[99]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[99])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_98 (
      .Q(out_o[98]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[98])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_97 (
      .Q(out_o[97]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[97])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_96 (
      .Q(out_o[96]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[96])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_95 (
      .Q(out_o[95]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[95])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_94 (
      .Q(out_o[94]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[94])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_93 (
      .Q(out_o[93]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[93])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_92 (
      .Q(out_o[92]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[92])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_91 (
      .Q(out_o[91]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[91])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_90 (
      .Q(out_o[90]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[90])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_89 (
      .Q(out_o[89]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[89])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_88 (
      .Q(out_o[88]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[88])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_87 (
      .Q(out_o[87]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[87])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_86 (
      .Q(out_o[86]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[86])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_85 (
      .Q(out_o[85]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[85])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_84 (
      .Q(out_o[84]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[84])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_83 (
      .Q(out_o[83]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[83])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_82 (
      .Q(out_o[82]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[82])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_81 (
      .Q(out_o[81]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[81])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_80 (
      .Q(out_o[80]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[80])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_79 (
      .Q(out_o[79]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[79])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_78 (
      .Q(out_o[78]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[78])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_77 (
      .Q(out_o[77]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[77])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_76 (
      .Q(out_o[76]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[76])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_75 (
      .Q(out_o[75]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[75])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_74 (
      .Q(out_o[74]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[74])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_73 (
      .Q(out_o[73]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[73])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_72 (
      .Q(out_o[72]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[72])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_71 (
      .Q(out_o[71]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[71])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_70 (
      .Q(out_o[70]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[70])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_69 (
      .Q(out_o[69]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[69])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_68 (
      .Q(out_o[68]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[68])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_67 (
      .Q(out_o[67]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[67])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_66 (
      .Q(out_o[66]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[66])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_65 (
      .Q(out_o[65]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[65])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_64 (
      .Q(out_o[64]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[64])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_63 (
      .Q(out_o[63]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[63])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_62 (
      .Q(out_o[62]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[62])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_61 (
      .Q(out_o[61]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[61])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_60 (
      .Q(out_o[60]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[60])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_59 (
      .Q(out_o[59]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[59])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_58 (
      .Q(out_o[58]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[58])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_57 (
      .Q(out_o[57]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[57])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_56 (
      .Q(out_o[56]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[56])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_55 (
      .Q(out_o[55]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[55])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_54 (
      .Q(out_o[54]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[54])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_53 (
      .Q(out_o[53]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[53])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_52 (
      .Q(out_o[52]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[52])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_51 (
      .Q(out_o[51]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[51])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_50 (
      .Q(out_o[50]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[50])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_49 (
      .Q(out_o[49]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[49])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_48 (
      .Q(out_o[48]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[48])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_47 (
      .Q(out_o[47]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[47])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_46 (
      .Q(out_o[46]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[46])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_45 (
      .Q(out_o[45]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[45])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_44 (
      .Q(out_o[44]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[44])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_43 (
      .Q(out_o[43]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[43])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_42 (
      .Q(out_o[42]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[42])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_41 (
      .Q(out_o[41]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[41])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_40 (
      .Q(out_o[40]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[40])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_39 (
      .Q(out_o[39]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[39])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_38 (
      .Q(out_o[38]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[38])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_37 (
      .Q(out_o[37]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[37])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_36 (
      .Q(out_o[36]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[36])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_35 (
      .Q(out_o[35]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[35])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_34 (
      .Q(out_o[34]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[34])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_33 (
      .Q(out_o[33]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[33])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_32 (
      .Q(out_o[32]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[32])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_31 (
      .Q(out_o[31]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[31])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_30 (
      .Q(out_o[30]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[30])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_29 (
      .Q(out_o[29]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[29])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_28 (
      .Q(out_o[28]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[28])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_27 (
      .Q(out_o[27]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[27])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_26 (
      .Q(out_o[26]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[26])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_25 (
      .Q(out_o[25]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[25])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_24 (
      .Q(out_o[24]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[24])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_23 (
      .Q(out_o[23]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[23])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_22 (
      .Q(out_o[22]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[22])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_21 (
      .Q(out_o[21]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[21])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_20 (
      .Q(out_o[20]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[20])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_19 (
      .Q(out_o[19]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[19])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_18 (
      .Q(out_o[18]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[18])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_17 (
      .Q(out_o[17]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[17])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_16 (
      .Q(out_o[16]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[16])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_15 (
      .Q(out_o[15]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[15])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_14 (
      .Q(out_o[14]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[14])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_13 (
      .Q(out_o[13]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[13])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_12 (
      .Q(out_o[12]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[12])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_11 (
      .Q(out_o[11]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[11])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_10 (
      .Q(out_o[10]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[10])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_9 (
      .Q(out_o[9]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[9])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_8 (
      .Q(out_o[8]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[8])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_7 (
      .Q(out_o[7]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[7])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_6 (
      .Q(out_o[6]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[6])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_5 (
      .Q(out_o[5]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[5])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_4 (
      .Q(out_o[4]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[4])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_3 (
      .Q(out_o[3]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[3])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_2 (
      .Q(out_o[2]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[2])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_1 (
      .Q(out_o[1]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[1])       // Data input
   );
       FDE #(
      .INIT(1'b0) // Initial value of register (1'b0 or 1'b1)
   ) out_o_0 (
      .Q(out_o[0]),      // Data output
      .C(clk_i),      // Clock input
      .CE(ce_i),    // Clock enable input
      .D(out[0])       // Data input
   );

endmodule

`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 05/17/2021 05:34:13 AM
// Design Name: 
// Module Name: mux_2i1o_512b
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module mux_2i1o_512b(
    input sel_i,
    input  [511:0] in_0_i,
    input  [511:0] in_1_i,

    output [511:0] out
    );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_511(.O(out[511]),     // LUT general output
                .I0(in_0_i[511]), // LUT input
                .I1(in_1_i[511]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_510(.O(out[510]),     // LUT general output
                .I0(in_0_i[510]), // LUT input
                .I1(in_1_i[510]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_509(.O(out[509]),     // LUT general output
                .I0(in_0_i[509]), // LUT input
                .I1(in_1_i[509]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_508(.O(out[508]),     // LUT general output
                .I0(in_0_i[508]), // LUT input
                .I1(in_1_i[508]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_507(.O(out[507]),     // LUT general output
                .I0(in_0_i[507]), // LUT input
                .I1(in_1_i[507]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_506(.O(out[506]),     // LUT general output
                .I0(in_0_i[506]), // LUT input
                .I1(in_1_i[506]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_505(.O(out[505]),     // LUT general output
                .I0(in_0_i[505]), // LUT input
                .I1(in_1_i[505]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_504(.O(out[504]),     // LUT general output
                .I0(in_0_i[504]), // LUT input
                .I1(in_1_i[504]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_503(.O(out[503]),     // LUT general output
                .I0(in_0_i[503]), // LUT input
                .I1(in_1_i[503]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_502(.O(out[502]),     // LUT general output
                .I0(in_0_i[502]), // LUT input
                .I1(in_1_i[502]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_501(.O(out[501]),     // LUT general output
                .I0(in_0_i[501]), // LUT input
                .I1(in_1_i[501]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_500(.O(out[500]),     // LUT general output
                .I0(in_0_i[500]), // LUT input
                .I1(in_1_i[500]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_499(.O(out[499]),     // LUT general output
                .I0(in_0_i[499]), // LUT input
                .I1(in_1_i[499]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_498(.O(out[498]),     // LUT general output
                .I0(in_0_i[498]), // LUT input
                .I1(in_1_i[498]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_497(.O(out[497]),     // LUT general output
                .I0(in_0_i[497]), // LUT input
                .I1(in_1_i[497]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_496(.O(out[496]),     // LUT general output
                .I0(in_0_i[496]), // LUT input
                .I1(in_1_i[496]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_495(.O(out[495]),     // LUT general output
                .I0(in_0_i[495]), // LUT input
                .I1(in_1_i[495]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_494(.O(out[494]),     // LUT general output
                .I0(in_0_i[494]), // LUT input
                .I1(in_1_i[494]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_493(.O(out[493]),     // LUT general output
                .I0(in_0_i[493]), // LUT input
                .I1(in_1_i[493]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_492(.O(out[492]),     // LUT general output
                .I0(in_0_i[492]), // LUT input
                .I1(in_1_i[492]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_491(.O(out[491]),     // LUT general output
                .I0(in_0_i[491]), // LUT input
                .I1(in_1_i[491]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_490(.O(out[490]),     // LUT general output
                .I0(in_0_i[490]), // LUT input
                .I1(in_1_i[490]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_489(.O(out[489]),     // LUT general output
                .I0(in_0_i[489]), // LUT input
                .I1(in_1_i[489]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_488(.O(out[488]),     // LUT general output
                .I0(in_0_i[488]), // LUT input
                .I1(in_1_i[488]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_487(.O(out[487]),     // LUT general output
                .I0(in_0_i[487]), // LUT input
                .I1(in_1_i[487]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_486(.O(out[486]),     // LUT general output
                .I0(in_0_i[486]), // LUT input
                .I1(in_1_i[486]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_485(.O(out[485]),     // LUT general output
                .I0(in_0_i[485]), // LUT input
                .I1(in_1_i[485]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_484(.O(out[484]),     // LUT general output
                .I0(in_0_i[484]), // LUT input
                .I1(in_1_i[484]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_483(.O(out[483]),     // LUT general output
                .I0(in_0_i[483]), // LUT input
                .I1(in_1_i[483]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_482(.O(out[482]),     // LUT general output
                .I0(in_0_i[482]), // LUT input
                .I1(in_1_i[482]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_481(.O(out[481]),     // LUT general output
                .I0(in_0_i[481]), // LUT input
                .I1(in_1_i[481]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_480(.O(out[480]),     // LUT general output
                .I0(in_0_i[480]), // LUT input
                .I1(in_1_i[480]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_479(.O(out[479]),     // LUT general output
                .I0(in_0_i[479]), // LUT input
                .I1(in_1_i[479]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_478(.O(out[478]),     // LUT general output
                .I0(in_0_i[478]), // LUT input
                .I1(in_1_i[478]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_477(.O(out[477]),     // LUT general output
                .I0(in_0_i[477]), // LUT input
                .I1(in_1_i[477]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_476(.O(out[476]),     // LUT general output
                .I0(in_0_i[476]), // LUT input
                .I1(in_1_i[476]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_475(.O(out[475]),     // LUT general output
                .I0(in_0_i[475]), // LUT input
                .I1(in_1_i[475]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_474(.O(out[474]),     // LUT general output
                .I0(in_0_i[474]), // LUT input
                .I1(in_1_i[474]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_473(.O(out[473]),     // LUT general output
                .I0(in_0_i[473]), // LUT input
                .I1(in_1_i[473]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_472(.O(out[472]),     // LUT general output
                .I0(in_0_i[472]), // LUT input
                .I1(in_1_i[472]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_471(.O(out[471]),     // LUT general output
                .I0(in_0_i[471]), // LUT input
                .I1(in_1_i[471]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_470(.O(out[470]),     // LUT general output
                .I0(in_0_i[470]), // LUT input
                .I1(in_1_i[470]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_469(.O(out[469]),     // LUT general output
                .I0(in_0_i[469]), // LUT input
                .I1(in_1_i[469]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_468(.O(out[468]),     // LUT general output
                .I0(in_0_i[468]), // LUT input
                .I1(in_1_i[468]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_467(.O(out[467]),     // LUT general output
                .I0(in_0_i[467]), // LUT input
                .I1(in_1_i[467]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_466(.O(out[466]),     // LUT general output
                .I0(in_0_i[466]), // LUT input
                .I1(in_1_i[466]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_465(.O(out[465]),     // LUT general output
                .I0(in_0_i[465]), // LUT input
                .I1(in_1_i[465]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_464(.O(out[464]),     // LUT general output
                .I0(in_0_i[464]), // LUT input
                .I1(in_1_i[464]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_463(.O(out[463]),     // LUT general output
                .I0(in_0_i[463]), // LUT input
                .I1(in_1_i[463]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_462(.O(out[462]),     // LUT general output
                .I0(in_0_i[462]), // LUT input
                .I1(in_1_i[462]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_461(.O(out[461]),     // LUT general output
                .I0(in_0_i[461]), // LUT input
                .I1(in_1_i[461]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_460(.O(out[460]),     // LUT general output
                .I0(in_0_i[460]), // LUT input
                .I1(in_1_i[460]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_459(.O(out[459]),     // LUT general output
                .I0(in_0_i[459]), // LUT input
                .I1(in_1_i[459]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_458(.O(out[458]),     // LUT general output
                .I0(in_0_i[458]), // LUT input
                .I1(in_1_i[458]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_457(.O(out[457]),     // LUT general output
                .I0(in_0_i[457]), // LUT input
                .I1(in_1_i[457]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_456(.O(out[456]),     // LUT general output
                .I0(in_0_i[456]), // LUT input
                .I1(in_1_i[456]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_455(.O(out[455]),     // LUT general output
                .I0(in_0_i[455]), // LUT input
                .I1(in_1_i[455]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_454(.O(out[454]),     // LUT general output
                .I0(in_0_i[454]), // LUT input
                .I1(in_1_i[454]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_453(.O(out[453]),     // LUT general output
                .I0(in_0_i[453]), // LUT input
                .I1(in_1_i[453]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_452(.O(out[452]),     // LUT general output
                .I0(in_0_i[452]), // LUT input
                .I1(in_1_i[452]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_451(.O(out[451]),     // LUT general output
                .I0(in_0_i[451]), // LUT input
                .I1(in_1_i[451]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_450(.O(out[450]),     // LUT general output
                .I0(in_0_i[450]), // LUT input
                .I1(in_1_i[450]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_449(.O(out[449]),     // LUT general output
                .I0(in_0_i[449]), // LUT input
                .I1(in_1_i[449]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_448(.O(out[448]),     // LUT general output
                .I0(in_0_i[448]), // LUT input
                .I1(in_1_i[448]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_447(.O(out[447]),     // LUT general output
                .I0(in_0_i[447]), // LUT input
                .I1(in_1_i[447]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_446(.O(out[446]),     // LUT general output
                .I0(in_0_i[446]), // LUT input
                .I1(in_1_i[446]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_445(.O(out[445]),     // LUT general output
                .I0(in_0_i[445]), // LUT input
                .I1(in_1_i[445]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_444(.O(out[444]),     // LUT general output
                .I0(in_0_i[444]), // LUT input
                .I1(in_1_i[444]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_443(.O(out[443]),     // LUT general output
                .I0(in_0_i[443]), // LUT input
                .I1(in_1_i[443]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_442(.O(out[442]),     // LUT general output
                .I0(in_0_i[442]), // LUT input
                .I1(in_1_i[442]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_441(.O(out[441]),     // LUT general output
                .I0(in_0_i[441]), // LUT input
                .I1(in_1_i[441]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_440(.O(out[440]),     // LUT general output
                .I0(in_0_i[440]), // LUT input
                .I1(in_1_i[440]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_439(.O(out[439]),     // LUT general output
                .I0(in_0_i[439]), // LUT input
                .I1(in_1_i[439]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_438(.O(out[438]),     // LUT general output
                .I0(in_0_i[438]), // LUT input
                .I1(in_1_i[438]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_437(.O(out[437]),     // LUT general output
                .I0(in_0_i[437]), // LUT input
                .I1(in_1_i[437]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_436(.O(out[436]),     // LUT general output
                .I0(in_0_i[436]), // LUT input
                .I1(in_1_i[436]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_435(.O(out[435]),     // LUT general output
                .I0(in_0_i[435]), // LUT input
                .I1(in_1_i[435]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_434(.O(out[434]),     // LUT general output
                .I0(in_0_i[434]), // LUT input
                .I1(in_1_i[434]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_433(.O(out[433]),     // LUT general output
                .I0(in_0_i[433]), // LUT input
                .I1(in_1_i[433]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_432(.O(out[432]),     // LUT general output
                .I0(in_0_i[432]), // LUT input
                .I1(in_1_i[432]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_431(.O(out[431]),     // LUT general output
                .I0(in_0_i[431]), // LUT input
                .I1(in_1_i[431]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_430(.O(out[430]),     // LUT general output
                .I0(in_0_i[430]), // LUT input
                .I1(in_1_i[430]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_429(.O(out[429]),     // LUT general output
                .I0(in_0_i[429]), // LUT input
                .I1(in_1_i[429]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_428(.O(out[428]),     // LUT general output
                .I0(in_0_i[428]), // LUT input
                .I1(in_1_i[428]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_427(.O(out[427]),     // LUT general output
                .I0(in_0_i[427]), // LUT input
                .I1(in_1_i[427]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_426(.O(out[426]),     // LUT general output
                .I0(in_0_i[426]), // LUT input
                .I1(in_1_i[426]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_425(.O(out[425]),     // LUT general output
                .I0(in_0_i[425]), // LUT input
                .I1(in_1_i[425]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_424(.O(out[424]),     // LUT general output
                .I0(in_0_i[424]), // LUT input
                .I1(in_1_i[424]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_423(.O(out[423]),     // LUT general output
                .I0(in_0_i[423]), // LUT input
                .I1(in_1_i[423]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_422(.O(out[422]),     // LUT general output
                .I0(in_0_i[422]), // LUT input
                .I1(in_1_i[422]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_421(.O(out[421]),     // LUT general output
                .I0(in_0_i[421]), // LUT input
                .I1(in_1_i[421]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_420(.O(out[420]),     // LUT general output
                .I0(in_0_i[420]), // LUT input
                .I1(in_1_i[420]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_419(.O(out[419]),     // LUT general output
                .I0(in_0_i[419]), // LUT input
                .I1(in_1_i[419]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_418(.O(out[418]),     // LUT general output
                .I0(in_0_i[418]), // LUT input
                .I1(in_1_i[418]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_417(.O(out[417]),     // LUT general output
                .I0(in_0_i[417]), // LUT input
                .I1(in_1_i[417]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_416(.O(out[416]),     // LUT general output
                .I0(in_0_i[416]), // LUT input
                .I1(in_1_i[416]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_415(.O(out[415]),     // LUT general output
                .I0(in_0_i[415]), // LUT input
                .I1(in_1_i[415]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_414(.O(out[414]),     // LUT general output
                .I0(in_0_i[414]), // LUT input
                .I1(in_1_i[414]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_413(.O(out[413]),     // LUT general output
                .I0(in_0_i[413]), // LUT input
                .I1(in_1_i[413]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_412(.O(out[412]),     // LUT general output
                .I0(in_0_i[412]), // LUT input
                .I1(in_1_i[412]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_411(.O(out[411]),     // LUT general output
                .I0(in_0_i[411]), // LUT input
                .I1(in_1_i[411]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_410(.O(out[410]),     // LUT general output
                .I0(in_0_i[410]), // LUT input
                .I1(in_1_i[410]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_409(.O(out[409]),     // LUT general output
                .I0(in_0_i[409]), // LUT input
                .I1(in_1_i[409]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_408(.O(out[408]),     // LUT general output
                .I0(in_0_i[408]), // LUT input
                .I1(in_1_i[408]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_407(.O(out[407]),     // LUT general output
                .I0(in_0_i[407]), // LUT input
                .I1(in_1_i[407]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_406(.O(out[406]),     // LUT general output
                .I0(in_0_i[406]), // LUT input
                .I1(in_1_i[406]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_405(.O(out[405]),     // LUT general output
                .I0(in_0_i[405]), // LUT input
                .I1(in_1_i[405]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_404(.O(out[404]),     // LUT general output
                .I0(in_0_i[404]), // LUT input
                .I1(in_1_i[404]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_403(.O(out[403]),     // LUT general output
                .I0(in_0_i[403]), // LUT input
                .I1(in_1_i[403]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_402(.O(out[402]),     // LUT general output
                .I0(in_0_i[402]), // LUT input
                .I1(in_1_i[402]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_401(.O(out[401]),     // LUT general output
                .I0(in_0_i[401]), // LUT input
                .I1(in_1_i[401]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_400(.O(out[400]),     // LUT general output
                .I0(in_0_i[400]), // LUT input
                .I1(in_1_i[400]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_399(.O(out[399]),     // LUT general output
                .I0(in_0_i[399]), // LUT input
                .I1(in_1_i[399]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_398(.O(out[398]),     // LUT general output
                .I0(in_0_i[398]), // LUT input
                .I1(in_1_i[398]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_397(.O(out[397]),     // LUT general output
                .I0(in_0_i[397]), // LUT input
                .I1(in_1_i[397]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_396(.O(out[396]),     // LUT general output
                .I0(in_0_i[396]), // LUT input
                .I1(in_1_i[396]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_395(.O(out[395]),     // LUT general output
                .I0(in_0_i[395]), // LUT input
                .I1(in_1_i[395]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_394(.O(out[394]),     // LUT general output
                .I0(in_0_i[394]), // LUT input
                .I1(in_1_i[394]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_393(.O(out[393]),     // LUT general output
                .I0(in_0_i[393]), // LUT input
                .I1(in_1_i[393]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_392(.O(out[392]),     // LUT general output
                .I0(in_0_i[392]), // LUT input
                .I1(in_1_i[392]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_391(.O(out[391]),     // LUT general output
                .I0(in_0_i[391]), // LUT input
                .I1(in_1_i[391]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_390(.O(out[390]),     // LUT general output
                .I0(in_0_i[390]), // LUT input
                .I1(in_1_i[390]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_389(.O(out[389]),     // LUT general output
                .I0(in_0_i[389]), // LUT input
                .I1(in_1_i[389]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_388(.O(out[388]),     // LUT general output
                .I0(in_0_i[388]), // LUT input
                .I1(in_1_i[388]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_387(.O(out[387]),     // LUT general output
                .I0(in_0_i[387]), // LUT input
                .I1(in_1_i[387]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_386(.O(out[386]),     // LUT general output
                .I0(in_0_i[386]), // LUT input
                .I1(in_1_i[386]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_385(.O(out[385]),     // LUT general output
                .I0(in_0_i[385]), // LUT input
                .I1(in_1_i[385]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_384(.O(out[384]),     // LUT general output
                .I0(in_0_i[384]), // LUT input
                .I1(in_1_i[384]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_383(.O(out[383]),     // LUT general output
                .I0(in_0_i[383]), // LUT input
                .I1(in_1_i[383]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_382(.O(out[382]),     // LUT general output
                .I0(in_0_i[382]), // LUT input
                .I1(in_1_i[382]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_381(.O(out[381]),     // LUT general output
                .I0(in_0_i[381]), // LUT input
                .I1(in_1_i[381]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_380(.O(out[380]),     // LUT general output
                .I0(in_0_i[380]), // LUT input
                .I1(in_1_i[380]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_379(.O(out[379]),     // LUT general output
                .I0(in_0_i[379]), // LUT input
                .I1(in_1_i[379]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_378(.O(out[378]),     // LUT general output
                .I0(in_0_i[378]), // LUT input
                .I1(in_1_i[378]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_377(.O(out[377]),     // LUT general output
                .I0(in_0_i[377]), // LUT input
                .I1(in_1_i[377]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_376(.O(out[376]),     // LUT general output
                .I0(in_0_i[376]), // LUT input
                .I1(in_1_i[376]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_375(.O(out[375]),     // LUT general output
                .I0(in_0_i[375]), // LUT input
                .I1(in_1_i[375]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_374(.O(out[374]),     // LUT general output
                .I0(in_0_i[374]), // LUT input
                .I1(in_1_i[374]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_373(.O(out[373]),     // LUT general output
                .I0(in_0_i[373]), // LUT input
                .I1(in_1_i[373]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_372(.O(out[372]),     // LUT general output
                .I0(in_0_i[372]), // LUT input
                .I1(in_1_i[372]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_371(.O(out[371]),     // LUT general output
                .I0(in_0_i[371]), // LUT input
                .I1(in_1_i[371]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_370(.O(out[370]),     // LUT general output
                .I0(in_0_i[370]), // LUT input
                .I1(in_1_i[370]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_369(.O(out[369]),     // LUT general output
                .I0(in_0_i[369]), // LUT input
                .I1(in_1_i[369]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_368(.O(out[368]),     // LUT general output
                .I0(in_0_i[368]), // LUT input
                .I1(in_1_i[368]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_367(.O(out[367]),     // LUT general output
                .I0(in_0_i[367]), // LUT input
                .I1(in_1_i[367]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_366(.O(out[366]),     // LUT general output
                .I0(in_0_i[366]), // LUT input
                .I1(in_1_i[366]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_365(.O(out[365]),     // LUT general output
                .I0(in_0_i[365]), // LUT input
                .I1(in_1_i[365]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_364(.O(out[364]),     // LUT general output
                .I0(in_0_i[364]), // LUT input
                .I1(in_1_i[364]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_363(.O(out[363]),     // LUT general output
                .I0(in_0_i[363]), // LUT input
                .I1(in_1_i[363]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_362(.O(out[362]),     // LUT general output
                .I0(in_0_i[362]), // LUT input
                .I1(in_1_i[362]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_361(.O(out[361]),     // LUT general output
                .I0(in_0_i[361]), // LUT input
                .I1(in_1_i[361]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_360(.O(out[360]),     // LUT general output
                .I0(in_0_i[360]), // LUT input
                .I1(in_1_i[360]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_359(.O(out[359]),     // LUT general output
                .I0(in_0_i[359]), // LUT input
                .I1(in_1_i[359]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_358(.O(out[358]),     // LUT general output
                .I0(in_0_i[358]), // LUT input
                .I1(in_1_i[358]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_357(.O(out[357]),     // LUT general output
                .I0(in_0_i[357]), // LUT input
                .I1(in_1_i[357]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_356(.O(out[356]),     // LUT general output
                .I0(in_0_i[356]), // LUT input
                .I1(in_1_i[356]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_355(.O(out[355]),     // LUT general output
                .I0(in_0_i[355]), // LUT input
                .I1(in_1_i[355]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_354(.O(out[354]),     // LUT general output
                .I0(in_0_i[354]), // LUT input
                .I1(in_1_i[354]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_353(.O(out[353]),     // LUT general output
                .I0(in_0_i[353]), // LUT input
                .I1(in_1_i[353]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_352(.O(out[352]),     // LUT general output
                .I0(in_0_i[352]), // LUT input
                .I1(in_1_i[352]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_351(.O(out[351]),     // LUT general output
                .I0(in_0_i[351]), // LUT input
                .I1(in_1_i[351]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_350(.O(out[350]),     // LUT general output
                .I0(in_0_i[350]), // LUT input
                .I1(in_1_i[350]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_349(.O(out[349]),     // LUT general output
                .I0(in_0_i[349]), // LUT input
                .I1(in_1_i[349]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_348(.O(out[348]),     // LUT general output
                .I0(in_0_i[348]), // LUT input
                .I1(in_1_i[348]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_347(.O(out[347]),     // LUT general output
                .I0(in_0_i[347]), // LUT input
                .I1(in_1_i[347]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_346(.O(out[346]),     // LUT general output
                .I0(in_0_i[346]), // LUT input
                .I1(in_1_i[346]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_345(.O(out[345]),     // LUT general output
                .I0(in_0_i[345]), // LUT input
                .I1(in_1_i[345]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_344(.O(out[344]),     // LUT general output
                .I0(in_0_i[344]), // LUT input
                .I1(in_1_i[344]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_343(.O(out[343]),     // LUT general output
                .I0(in_0_i[343]), // LUT input
                .I1(in_1_i[343]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_342(.O(out[342]),     // LUT general output
                .I0(in_0_i[342]), // LUT input
                .I1(in_1_i[342]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_341(.O(out[341]),     // LUT general output
                .I0(in_0_i[341]), // LUT input
                .I1(in_1_i[341]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_340(.O(out[340]),     // LUT general output
                .I0(in_0_i[340]), // LUT input
                .I1(in_1_i[340]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_339(.O(out[339]),     // LUT general output
                .I0(in_0_i[339]), // LUT input
                .I1(in_1_i[339]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_338(.O(out[338]),     // LUT general output
                .I0(in_0_i[338]), // LUT input
                .I1(in_1_i[338]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_337(.O(out[337]),     // LUT general output
                .I0(in_0_i[337]), // LUT input
                .I1(in_1_i[337]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_336(.O(out[336]),     // LUT general output
                .I0(in_0_i[336]), // LUT input
                .I1(in_1_i[336]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_335(.O(out[335]),     // LUT general output
                .I0(in_0_i[335]), // LUT input
                .I1(in_1_i[335]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_334(.O(out[334]),     // LUT general output
                .I0(in_0_i[334]), // LUT input
                .I1(in_1_i[334]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_333(.O(out[333]),     // LUT general output
                .I0(in_0_i[333]), // LUT input
                .I1(in_1_i[333]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_332(.O(out[332]),     // LUT general output
                .I0(in_0_i[332]), // LUT input
                .I1(in_1_i[332]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_331(.O(out[331]),     // LUT general output
                .I0(in_0_i[331]), // LUT input
                .I1(in_1_i[331]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_330(.O(out[330]),     // LUT general output
                .I0(in_0_i[330]), // LUT input
                .I1(in_1_i[330]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_329(.O(out[329]),     // LUT general output
                .I0(in_0_i[329]), // LUT input
                .I1(in_1_i[329]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_328(.O(out[328]),     // LUT general output
                .I0(in_0_i[328]), // LUT input
                .I1(in_1_i[328]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_327(.O(out[327]),     // LUT general output
                .I0(in_0_i[327]), // LUT input
                .I1(in_1_i[327]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_326(.O(out[326]),     // LUT general output
                .I0(in_0_i[326]), // LUT input
                .I1(in_1_i[326]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_325(.O(out[325]),     // LUT general output
                .I0(in_0_i[325]), // LUT input
                .I1(in_1_i[325]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_324(.O(out[324]),     // LUT general output
                .I0(in_0_i[324]), // LUT input
                .I1(in_1_i[324]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_323(.O(out[323]),     // LUT general output
                .I0(in_0_i[323]), // LUT input
                .I1(in_1_i[323]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_322(.O(out[322]),     // LUT general output
                .I0(in_0_i[322]), // LUT input
                .I1(in_1_i[322]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_321(.O(out[321]),     // LUT general output
                .I0(in_0_i[321]), // LUT input
                .I1(in_1_i[321]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_320(.O(out[320]),     // LUT general output
                .I0(in_0_i[320]), // LUT input
                .I1(in_1_i[320]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_319(.O(out[319]),     // LUT general output
                .I0(in_0_i[319]), // LUT input
                .I1(in_1_i[319]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_318(.O(out[318]),     // LUT general output
                .I0(in_0_i[318]), // LUT input
                .I1(in_1_i[318]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_317(.O(out[317]),     // LUT general output
                .I0(in_0_i[317]), // LUT input
                .I1(in_1_i[317]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_316(.O(out[316]),     // LUT general output
                .I0(in_0_i[316]), // LUT input
                .I1(in_1_i[316]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_315(.O(out[315]),     // LUT general output
                .I0(in_0_i[315]), // LUT input
                .I1(in_1_i[315]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_314(.O(out[314]),     // LUT general output
                .I0(in_0_i[314]), // LUT input
                .I1(in_1_i[314]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_313(.O(out[313]),     // LUT general output
                .I0(in_0_i[313]), // LUT input
                .I1(in_1_i[313]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_312(.O(out[312]),     // LUT general output
                .I0(in_0_i[312]), // LUT input
                .I1(in_1_i[312]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_311(.O(out[311]),     // LUT general output
                .I0(in_0_i[311]), // LUT input
                .I1(in_1_i[311]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_310(.O(out[310]),     // LUT general output
                .I0(in_0_i[310]), // LUT input
                .I1(in_1_i[310]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_309(.O(out[309]),     // LUT general output
                .I0(in_0_i[309]), // LUT input
                .I1(in_1_i[309]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_308(.O(out[308]),     // LUT general output
                .I0(in_0_i[308]), // LUT input
                .I1(in_1_i[308]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_307(.O(out[307]),     // LUT general output
                .I0(in_0_i[307]), // LUT input
                .I1(in_1_i[307]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_306(.O(out[306]),     // LUT general output
                .I0(in_0_i[306]), // LUT input
                .I1(in_1_i[306]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_305(.O(out[305]),     // LUT general output
                .I0(in_0_i[305]), // LUT input
                .I1(in_1_i[305]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_304(.O(out[304]),     // LUT general output
                .I0(in_0_i[304]), // LUT input
                .I1(in_1_i[304]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_303(.O(out[303]),     // LUT general output
                .I0(in_0_i[303]), // LUT input
                .I1(in_1_i[303]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_302(.O(out[302]),     // LUT general output
                .I0(in_0_i[302]), // LUT input
                .I1(in_1_i[302]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_301(.O(out[301]),     // LUT general output
                .I0(in_0_i[301]), // LUT input
                .I1(in_1_i[301]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_300(.O(out[300]),     // LUT general output
                .I0(in_0_i[300]), // LUT input
                .I1(in_1_i[300]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_299(.O(out[299]),     // LUT general output
                .I0(in_0_i[299]), // LUT input
                .I1(in_1_i[299]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_298(.O(out[298]),     // LUT general output
                .I0(in_0_i[298]), // LUT input
                .I1(in_1_i[298]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_297(.O(out[297]),     // LUT general output
                .I0(in_0_i[297]), // LUT input
                .I1(in_1_i[297]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_296(.O(out[296]),     // LUT general output
                .I0(in_0_i[296]), // LUT input
                .I1(in_1_i[296]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_295(.O(out[295]),     // LUT general output
                .I0(in_0_i[295]), // LUT input
                .I1(in_1_i[295]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_294(.O(out[294]),     // LUT general output
                .I0(in_0_i[294]), // LUT input
                .I1(in_1_i[294]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_293(.O(out[293]),     // LUT general output
                .I0(in_0_i[293]), // LUT input
                .I1(in_1_i[293]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_292(.O(out[292]),     // LUT general output
                .I0(in_0_i[292]), // LUT input
                .I1(in_1_i[292]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_291(.O(out[291]),     // LUT general output
                .I0(in_0_i[291]), // LUT input
                .I1(in_1_i[291]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_290(.O(out[290]),     // LUT general output
                .I0(in_0_i[290]), // LUT input
                .I1(in_1_i[290]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_289(.O(out[289]),     // LUT general output
                .I0(in_0_i[289]), // LUT input
                .I1(in_1_i[289]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_288(.O(out[288]),     // LUT general output
                .I0(in_0_i[288]), // LUT input
                .I1(in_1_i[288]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_287(.O(out[287]),     // LUT general output
                .I0(in_0_i[287]), // LUT input
                .I1(in_1_i[287]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_286(.O(out[286]),     // LUT general output
                .I0(in_0_i[286]), // LUT input
                .I1(in_1_i[286]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_285(.O(out[285]),     // LUT general output
                .I0(in_0_i[285]), // LUT input
                .I1(in_1_i[285]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_284(.O(out[284]),     // LUT general output
                .I0(in_0_i[284]), // LUT input
                .I1(in_1_i[284]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_283(.O(out[283]),     // LUT general output
                .I0(in_0_i[283]), // LUT input
                .I1(in_1_i[283]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_282(.O(out[282]),     // LUT general output
                .I0(in_0_i[282]), // LUT input
                .I1(in_1_i[282]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_281(.O(out[281]),     // LUT general output
                .I0(in_0_i[281]), // LUT input
                .I1(in_1_i[281]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_280(.O(out[280]),     // LUT general output
                .I0(in_0_i[280]), // LUT input
                .I1(in_1_i[280]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_279(.O(out[279]),     // LUT general output
                .I0(in_0_i[279]), // LUT input
                .I1(in_1_i[279]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_278(.O(out[278]),     // LUT general output
                .I0(in_0_i[278]), // LUT input
                .I1(in_1_i[278]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_277(.O(out[277]),     // LUT general output
                .I0(in_0_i[277]), // LUT input
                .I1(in_1_i[277]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_276(.O(out[276]),     // LUT general output
                .I0(in_0_i[276]), // LUT input
                .I1(in_1_i[276]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_275(.O(out[275]),     // LUT general output
                .I0(in_0_i[275]), // LUT input
                .I1(in_1_i[275]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_274(.O(out[274]),     // LUT general output
                .I0(in_0_i[274]), // LUT input
                .I1(in_1_i[274]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_273(.O(out[273]),     // LUT general output
                .I0(in_0_i[273]), // LUT input
                .I1(in_1_i[273]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_272(.O(out[272]),     // LUT general output
                .I0(in_0_i[272]), // LUT input
                .I1(in_1_i[272]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_271(.O(out[271]),     // LUT general output
                .I0(in_0_i[271]), // LUT input
                .I1(in_1_i[271]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_270(.O(out[270]),     // LUT general output
                .I0(in_0_i[270]), // LUT input
                .I1(in_1_i[270]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_269(.O(out[269]),     // LUT general output
                .I0(in_0_i[269]), // LUT input
                .I1(in_1_i[269]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_268(.O(out[268]),     // LUT general output
                .I0(in_0_i[268]), // LUT input
                .I1(in_1_i[268]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_267(.O(out[267]),     // LUT general output
                .I0(in_0_i[267]), // LUT input
                .I1(in_1_i[267]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_266(.O(out[266]),     // LUT general output
                .I0(in_0_i[266]), // LUT input
                .I1(in_1_i[266]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_265(.O(out[265]),     // LUT general output
                .I0(in_0_i[265]), // LUT input
                .I1(in_1_i[265]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_264(.O(out[264]),     // LUT general output
                .I0(in_0_i[264]), // LUT input
                .I1(in_1_i[264]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_263(.O(out[263]),     // LUT general output
                .I0(in_0_i[263]), // LUT input
                .I1(in_1_i[263]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_262(.O(out[262]),     // LUT general output
                .I0(in_0_i[262]), // LUT input
                .I1(in_1_i[262]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_261(.O(out[261]),     // LUT general output
                .I0(in_0_i[261]), // LUT input
                .I1(in_1_i[261]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_260(.O(out[260]),     // LUT general output
                .I0(in_0_i[260]), // LUT input
                .I1(in_1_i[260]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_259(.O(out[259]),     // LUT general output
                .I0(in_0_i[259]), // LUT input
                .I1(in_1_i[259]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_258(.O(out[258]),     // LUT general output
                .I0(in_0_i[258]), // LUT input
                .I1(in_1_i[258]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_257(.O(out[257]),     // LUT general output
                .I0(in_0_i[257]), // LUT input
                .I1(in_1_i[257]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_256(.O(out[256]),     // LUT general output
                .I0(in_0_i[256]), // LUT input
                .I1(in_1_i[256]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_255(.O(out[255]),     // LUT general output
                .I0(in_0_i[255]), // LUT input
                .I1(in_1_i[255]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_254(.O(out[254]),     // LUT general output
                .I0(in_0_i[254]), // LUT input
                .I1(in_1_i[254]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_253(.O(out[253]),     // LUT general output
                .I0(in_0_i[253]), // LUT input
                .I1(in_1_i[253]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_252(.O(out[252]),     // LUT general output
                .I0(in_0_i[252]), // LUT input
                .I1(in_1_i[252]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_251(.O(out[251]),     // LUT general output
                .I0(in_0_i[251]), // LUT input
                .I1(in_1_i[251]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_250(.O(out[250]),     // LUT general output
                .I0(in_0_i[250]), // LUT input
                .I1(in_1_i[250]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_249(.O(out[249]),     // LUT general output
                .I0(in_0_i[249]), // LUT input
                .I1(in_1_i[249]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_248(.O(out[248]),     // LUT general output
                .I0(in_0_i[248]), // LUT input
                .I1(in_1_i[248]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_247(.O(out[247]),     // LUT general output
                .I0(in_0_i[247]), // LUT input
                .I1(in_1_i[247]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_246(.O(out[246]),     // LUT general output
                .I0(in_0_i[246]), // LUT input
                .I1(in_1_i[246]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_245(.O(out[245]),     // LUT general output
                .I0(in_0_i[245]), // LUT input
                .I1(in_1_i[245]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_244(.O(out[244]),     // LUT general output
                .I0(in_0_i[244]), // LUT input
                .I1(in_1_i[244]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_243(.O(out[243]),     // LUT general output
                .I0(in_0_i[243]), // LUT input
                .I1(in_1_i[243]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_242(.O(out[242]),     // LUT general output
                .I0(in_0_i[242]), // LUT input
                .I1(in_1_i[242]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_241(.O(out[241]),     // LUT general output
                .I0(in_0_i[241]), // LUT input
                .I1(in_1_i[241]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_240(.O(out[240]),     // LUT general output
                .I0(in_0_i[240]), // LUT input
                .I1(in_1_i[240]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_239(.O(out[239]),     // LUT general output
                .I0(in_0_i[239]), // LUT input
                .I1(in_1_i[239]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_238(.O(out[238]),     // LUT general output
                .I0(in_0_i[238]), // LUT input
                .I1(in_1_i[238]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_237(.O(out[237]),     // LUT general output
                .I0(in_0_i[237]), // LUT input
                .I1(in_1_i[237]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_236(.O(out[236]),     // LUT general output
                .I0(in_0_i[236]), // LUT input
                .I1(in_1_i[236]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_235(.O(out[235]),     // LUT general output
                .I0(in_0_i[235]), // LUT input
                .I1(in_1_i[235]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_234(.O(out[234]),     // LUT general output
                .I0(in_0_i[234]), // LUT input
                .I1(in_1_i[234]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_233(.O(out[233]),     // LUT general output
                .I0(in_0_i[233]), // LUT input
                .I1(in_1_i[233]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_232(.O(out[232]),     // LUT general output
                .I0(in_0_i[232]), // LUT input
                .I1(in_1_i[232]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_231(.O(out[231]),     // LUT general output
                .I0(in_0_i[231]), // LUT input
                .I1(in_1_i[231]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_230(.O(out[230]),     // LUT general output
                .I0(in_0_i[230]), // LUT input
                .I1(in_1_i[230]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_229(.O(out[229]),     // LUT general output
                .I0(in_0_i[229]), // LUT input
                .I1(in_1_i[229]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_228(.O(out[228]),     // LUT general output
                .I0(in_0_i[228]), // LUT input
                .I1(in_1_i[228]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_227(.O(out[227]),     // LUT general output
                .I0(in_0_i[227]), // LUT input
                .I1(in_1_i[227]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_226(.O(out[226]),     // LUT general output
                .I0(in_0_i[226]), // LUT input
                .I1(in_1_i[226]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_225(.O(out[225]),     // LUT general output
                .I0(in_0_i[225]), // LUT input
                .I1(in_1_i[225]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_224(.O(out[224]),     // LUT general output
                .I0(in_0_i[224]), // LUT input
                .I1(in_1_i[224]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_223(.O(out[223]),     // LUT general output
                .I0(in_0_i[223]), // LUT input
                .I1(in_1_i[223]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_222(.O(out[222]),     // LUT general output
                .I0(in_0_i[222]), // LUT input
                .I1(in_1_i[222]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_221(.O(out[221]),     // LUT general output
                .I0(in_0_i[221]), // LUT input
                .I1(in_1_i[221]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_220(.O(out[220]),     // LUT general output
                .I0(in_0_i[220]), // LUT input
                .I1(in_1_i[220]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_219(.O(out[219]),     // LUT general output
                .I0(in_0_i[219]), // LUT input
                .I1(in_1_i[219]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_218(.O(out[218]),     // LUT general output
                .I0(in_0_i[218]), // LUT input
                .I1(in_1_i[218]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_217(.O(out[217]),     // LUT general output
                .I0(in_0_i[217]), // LUT input
                .I1(in_1_i[217]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_216(.O(out[216]),     // LUT general output
                .I0(in_0_i[216]), // LUT input
                .I1(in_1_i[216]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_215(.O(out[215]),     // LUT general output
                .I0(in_0_i[215]), // LUT input
                .I1(in_1_i[215]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_214(.O(out[214]),     // LUT general output
                .I0(in_0_i[214]), // LUT input
                .I1(in_1_i[214]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_213(.O(out[213]),     // LUT general output
                .I0(in_0_i[213]), // LUT input
                .I1(in_1_i[213]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_212(.O(out[212]),     // LUT general output
                .I0(in_0_i[212]), // LUT input
                .I1(in_1_i[212]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_211(.O(out[211]),     // LUT general output
                .I0(in_0_i[211]), // LUT input
                .I1(in_1_i[211]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_210(.O(out[210]),     // LUT general output
                .I0(in_0_i[210]), // LUT input
                .I1(in_1_i[210]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_209(.O(out[209]),     // LUT general output
                .I0(in_0_i[209]), // LUT input
                .I1(in_1_i[209]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_208(.O(out[208]),     // LUT general output
                .I0(in_0_i[208]), // LUT input
                .I1(in_1_i[208]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_207(.O(out[207]),     // LUT general output
                .I0(in_0_i[207]), // LUT input
                .I1(in_1_i[207]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_206(.O(out[206]),     // LUT general output
                .I0(in_0_i[206]), // LUT input
                .I1(in_1_i[206]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_205(.O(out[205]),     // LUT general output
                .I0(in_0_i[205]), // LUT input
                .I1(in_1_i[205]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_204(.O(out[204]),     // LUT general output
                .I0(in_0_i[204]), // LUT input
                .I1(in_1_i[204]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_203(.O(out[203]),     // LUT general output
                .I0(in_0_i[203]), // LUT input
                .I1(in_1_i[203]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_202(.O(out[202]),     // LUT general output
                .I0(in_0_i[202]), // LUT input
                .I1(in_1_i[202]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_201(.O(out[201]),     // LUT general output
                .I0(in_0_i[201]), // LUT input
                .I1(in_1_i[201]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_200(.O(out[200]),     // LUT general output
                .I0(in_0_i[200]), // LUT input
                .I1(in_1_i[200]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_199(.O(out[199]),     // LUT general output
                .I0(in_0_i[199]), // LUT input
                .I1(in_1_i[199]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_198(.O(out[198]),     // LUT general output
                .I0(in_0_i[198]), // LUT input
                .I1(in_1_i[198]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_197(.O(out[197]),     // LUT general output
                .I0(in_0_i[197]), // LUT input
                .I1(in_1_i[197]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_196(.O(out[196]),     // LUT general output
                .I0(in_0_i[196]), // LUT input
                .I1(in_1_i[196]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_195(.O(out[195]),     // LUT general output
                .I0(in_0_i[195]), // LUT input
                .I1(in_1_i[195]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_194(.O(out[194]),     // LUT general output
                .I0(in_0_i[194]), // LUT input
                .I1(in_1_i[194]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_193(.O(out[193]),     // LUT general output
                .I0(in_0_i[193]), // LUT input
                .I1(in_1_i[193]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_192(.O(out[192]),     // LUT general output
                .I0(in_0_i[192]), // LUT input
                .I1(in_1_i[192]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_191(.O(out[191]),     // LUT general output
                .I0(in_0_i[191]), // LUT input
                .I1(in_1_i[191]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_190(.O(out[190]),     // LUT general output
                .I0(in_0_i[190]), // LUT input
                .I1(in_1_i[190]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_189(.O(out[189]),     // LUT general output
                .I0(in_0_i[189]), // LUT input
                .I1(in_1_i[189]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_188(.O(out[188]),     // LUT general output
                .I0(in_0_i[188]), // LUT input
                .I1(in_1_i[188]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_187(.O(out[187]),     // LUT general output
                .I0(in_0_i[187]), // LUT input
                .I1(in_1_i[187]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_186(.O(out[186]),     // LUT general output
                .I0(in_0_i[186]), // LUT input
                .I1(in_1_i[186]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_185(.O(out[185]),     // LUT general output
                .I0(in_0_i[185]), // LUT input
                .I1(in_1_i[185]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_184(.O(out[184]),     // LUT general output
                .I0(in_0_i[184]), // LUT input
                .I1(in_1_i[184]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_183(.O(out[183]),     // LUT general output
                .I0(in_0_i[183]), // LUT input
                .I1(in_1_i[183]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_182(.O(out[182]),     // LUT general output
                .I0(in_0_i[182]), // LUT input
                .I1(in_1_i[182]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_181(.O(out[181]),     // LUT general output
                .I0(in_0_i[181]), // LUT input
                .I1(in_1_i[181]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_180(.O(out[180]),     // LUT general output
                .I0(in_0_i[180]), // LUT input
                .I1(in_1_i[180]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_179(.O(out[179]),     // LUT general output
                .I0(in_0_i[179]), // LUT input
                .I1(in_1_i[179]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_178(.O(out[178]),     // LUT general output
                .I0(in_0_i[178]), // LUT input
                .I1(in_1_i[178]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_177(.O(out[177]),     // LUT general output
                .I0(in_0_i[177]), // LUT input
                .I1(in_1_i[177]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_176(.O(out[176]),     // LUT general output
                .I0(in_0_i[176]), // LUT input
                .I1(in_1_i[176]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_175(.O(out[175]),     // LUT general output
                .I0(in_0_i[175]), // LUT input
                .I1(in_1_i[175]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_174(.O(out[174]),     // LUT general output
                .I0(in_0_i[174]), // LUT input
                .I1(in_1_i[174]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_173(.O(out[173]),     // LUT general output
                .I0(in_0_i[173]), // LUT input
                .I1(in_1_i[173]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_172(.O(out[172]),     // LUT general output
                .I0(in_0_i[172]), // LUT input
                .I1(in_1_i[172]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_171(.O(out[171]),     // LUT general output
                .I0(in_0_i[171]), // LUT input
                .I1(in_1_i[171]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_170(.O(out[170]),     // LUT general output
                .I0(in_0_i[170]), // LUT input
                .I1(in_1_i[170]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_169(.O(out[169]),     // LUT general output
                .I0(in_0_i[169]), // LUT input
                .I1(in_1_i[169]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_168(.O(out[168]),     // LUT general output
                .I0(in_0_i[168]), // LUT input
                .I1(in_1_i[168]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_167(.O(out[167]),     // LUT general output
                .I0(in_0_i[167]), // LUT input
                .I1(in_1_i[167]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_166(.O(out[166]),     // LUT general output
                .I0(in_0_i[166]), // LUT input
                .I1(in_1_i[166]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_165(.O(out[165]),     // LUT general output
                .I0(in_0_i[165]), // LUT input
                .I1(in_1_i[165]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_164(.O(out[164]),     // LUT general output
                .I0(in_0_i[164]), // LUT input
                .I1(in_1_i[164]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_163(.O(out[163]),     // LUT general output
                .I0(in_0_i[163]), // LUT input
                .I1(in_1_i[163]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_162(.O(out[162]),     // LUT general output
                .I0(in_0_i[162]), // LUT input
                .I1(in_1_i[162]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_161(.O(out[161]),     // LUT general output
                .I0(in_0_i[161]), // LUT input
                .I1(in_1_i[161]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_160(.O(out[160]),     // LUT general output
                .I0(in_0_i[160]), // LUT input
                .I1(in_1_i[160]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_159(.O(out[159]),     // LUT general output
                .I0(in_0_i[159]), // LUT input
                .I1(in_1_i[159]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_158(.O(out[158]),     // LUT general output
                .I0(in_0_i[158]), // LUT input
                .I1(in_1_i[158]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_157(.O(out[157]),     // LUT general output
                .I0(in_0_i[157]), // LUT input
                .I1(in_1_i[157]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_156(.O(out[156]),     // LUT general output
                .I0(in_0_i[156]), // LUT input
                .I1(in_1_i[156]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_155(.O(out[155]),     // LUT general output
                .I0(in_0_i[155]), // LUT input
                .I1(in_1_i[155]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_154(.O(out[154]),     // LUT general output
                .I0(in_0_i[154]), // LUT input
                .I1(in_1_i[154]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_153(.O(out[153]),     // LUT general output
                .I0(in_0_i[153]), // LUT input
                .I1(in_1_i[153]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_152(.O(out[152]),     // LUT general output
                .I0(in_0_i[152]), // LUT input
                .I1(in_1_i[152]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_151(.O(out[151]),     // LUT general output
                .I0(in_0_i[151]), // LUT input
                .I1(in_1_i[151]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_150(.O(out[150]),     // LUT general output
                .I0(in_0_i[150]), // LUT input
                .I1(in_1_i[150]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_149(.O(out[149]),     // LUT general output
                .I0(in_0_i[149]), // LUT input
                .I1(in_1_i[149]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_148(.O(out[148]),     // LUT general output
                .I0(in_0_i[148]), // LUT input
                .I1(in_1_i[148]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_147(.O(out[147]),     // LUT general output
                .I0(in_0_i[147]), // LUT input
                .I1(in_1_i[147]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_146(.O(out[146]),     // LUT general output
                .I0(in_0_i[146]), // LUT input
                .I1(in_1_i[146]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_145(.O(out[145]),     // LUT general output
                .I0(in_0_i[145]), // LUT input
                .I1(in_1_i[145]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_144(.O(out[144]),     // LUT general output
                .I0(in_0_i[144]), // LUT input
                .I1(in_1_i[144]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_143(.O(out[143]),     // LUT general output
                .I0(in_0_i[143]), // LUT input
                .I1(in_1_i[143]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_142(.O(out[142]),     // LUT general output
                .I0(in_0_i[142]), // LUT input
                .I1(in_1_i[142]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_141(.O(out[141]),     // LUT general output
                .I0(in_0_i[141]), // LUT input
                .I1(in_1_i[141]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_140(.O(out[140]),     // LUT general output
                .I0(in_0_i[140]), // LUT input
                .I1(in_1_i[140]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_139(.O(out[139]),     // LUT general output
                .I0(in_0_i[139]), // LUT input
                .I1(in_1_i[139]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_138(.O(out[138]),     // LUT general output
                .I0(in_0_i[138]), // LUT input
                .I1(in_1_i[138]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_137(.O(out[137]),     // LUT general output
                .I0(in_0_i[137]), // LUT input
                .I1(in_1_i[137]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_136(.O(out[136]),     // LUT general output
                .I0(in_0_i[136]), // LUT input
                .I1(in_1_i[136]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_135(.O(out[135]),     // LUT general output
                .I0(in_0_i[135]), // LUT input
                .I1(in_1_i[135]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_134(.O(out[134]),     // LUT general output
                .I0(in_0_i[134]), // LUT input
                .I1(in_1_i[134]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_133(.O(out[133]),     // LUT general output
                .I0(in_0_i[133]), // LUT input
                .I1(in_1_i[133]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_132(.O(out[132]),     // LUT general output
                .I0(in_0_i[132]), // LUT input
                .I1(in_1_i[132]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_131(.O(out[131]),     // LUT general output
                .I0(in_0_i[131]), // LUT input
                .I1(in_1_i[131]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_130(.O(out[130]),     // LUT general output
                .I0(in_0_i[130]), // LUT input
                .I1(in_1_i[130]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_129(.O(out[129]),     // LUT general output
                .I0(in_0_i[129]), // LUT input
                .I1(in_1_i[129]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_128(.O(out[128]),     // LUT general output
                .I0(in_0_i[128]), // LUT input
                .I1(in_1_i[128]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_127(.O(out[127]),     // LUT general output
                .I0(in_0_i[127]), // LUT input
                .I1(in_1_i[127]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_126(.O(out[126]),     // LUT general output
                .I0(in_0_i[126]), // LUT input
                .I1(in_1_i[126]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_125(.O(out[125]),     // LUT general output
                .I0(in_0_i[125]), // LUT input
                .I1(in_1_i[125]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_124(.O(out[124]),     // LUT general output
                .I0(in_0_i[124]), // LUT input
                .I1(in_1_i[124]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_123(.O(out[123]),     // LUT general output
                .I0(in_0_i[123]), // LUT input
                .I1(in_1_i[123]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_122(.O(out[122]),     // LUT general output
                .I0(in_0_i[122]), // LUT input
                .I1(in_1_i[122]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_121(.O(out[121]),     // LUT general output
                .I0(in_0_i[121]), // LUT input
                .I1(in_1_i[121]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_120(.O(out[120]),     // LUT general output
                .I0(in_0_i[120]), // LUT input
                .I1(in_1_i[120]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_119(.O(out[119]),     // LUT general output
                .I0(in_0_i[119]), // LUT input
                .I1(in_1_i[119]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_118(.O(out[118]),     // LUT general output
                .I0(in_0_i[118]), // LUT input
                .I1(in_1_i[118]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_117(.O(out[117]),     // LUT general output
                .I0(in_0_i[117]), // LUT input
                .I1(in_1_i[117]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_116(.O(out[116]),     // LUT general output
                .I0(in_0_i[116]), // LUT input
                .I1(in_1_i[116]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_115(.O(out[115]),     // LUT general output
                .I0(in_0_i[115]), // LUT input
                .I1(in_1_i[115]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_114(.O(out[114]),     // LUT general output
                .I0(in_0_i[114]), // LUT input
                .I1(in_1_i[114]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_113(.O(out[113]),     // LUT general output
                .I0(in_0_i[113]), // LUT input
                .I1(in_1_i[113]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_112(.O(out[112]),     // LUT general output
                .I0(in_0_i[112]), // LUT input
                .I1(in_1_i[112]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_111(.O(out[111]),     // LUT general output
                .I0(in_0_i[111]), // LUT input
                .I1(in_1_i[111]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_110(.O(out[110]),     // LUT general output
                .I0(in_0_i[110]), // LUT input
                .I1(in_1_i[110]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_109(.O(out[109]),     // LUT general output
                .I0(in_0_i[109]), // LUT input
                .I1(in_1_i[109]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_108(.O(out[108]),     // LUT general output
                .I0(in_0_i[108]), // LUT input
                .I1(in_1_i[108]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_107(.O(out[107]),     // LUT general output
                .I0(in_0_i[107]), // LUT input
                .I1(in_1_i[107]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_106(.O(out[106]),     // LUT general output
                .I0(in_0_i[106]), // LUT input
                .I1(in_1_i[106]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_105(.O(out[105]),     // LUT general output
                .I0(in_0_i[105]), // LUT input
                .I1(in_1_i[105]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_104(.O(out[104]),     // LUT general output
                .I0(in_0_i[104]), // LUT input
                .I1(in_1_i[104]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_103(.O(out[103]),     // LUT general output
                .I0(in_0_i[103]), // LUT input
                .I1(in_1_i[103]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_102(.O(out[102]),     // LUT general output
                .I0(in_0_i[102]), // LUT input
                .I1(in_1_i[102]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_101(.O(out[101]),     // LUT general output
                .I0(in_0_i[101]), // LUT input
                .I1(in_1_i[101]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_100(.O(out[100]),     // LUT general output
                .I0(in_0_i[100]), // LUT input
                .I1(in_1_i[100]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_99(.O(out[99]),     // LUT general output
                .I0(in_0_i[99]), // LUT input
                .I1(in_1_i[99]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_98(.O(out[98]),     // LUT general output
                .I0(in_0_i[98]), // LUT input
                .I1(in_1_i[98]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_97(.O(out[97]),     // LUT general output
                .I0(in_0_i[97]), // LUT input
                .I1(in_1_i[97]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_96(.O(out[96]),     // LUT general output
                .I0(in_0_i[96]), // LUT input
                .I1(in_1_i[96]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_95(.O(out[95]),     // LUT general output
                .I0(in_0_i[95]), // LUT input
                .I1(in_1_i[95]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_94(.O(out[94]),     // LUT general output
                .I0(in_0_i[94]), // LUT input
                .I1(in_1_i[94]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_93(.O(out[93]),     // LUT general output
                .I0(in_0_i[93]), // LUT input
                .I1(in_1_i[93]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_92(.O(out[92]),     // LUT general output
                .I0(in_0_i[92]), // LUT input
                .I1(in_1_i[92]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_91(.O(out[91]),     // LUT general output
                .I0(in_0_i[91]), // LUT input
                .I1(in_1_i[91]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_90(.O(out[90]),     // LUT general output
                .I0(in_0_i[90]), // LUT input
                .I1(in_1_i[90]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_89(.O(out[89]),     // LUT general output
                .I0(in_0_i[89]), // LUT input
                .I1(in_1_i[89]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_88(.O(out[88]),     // LUT general output
                .I0(in_0_i[88]), // LUT input
                .I1(in_1_i[88]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_87(.O(out[87]),     // LUT general output
                .I0(in_0_i[87]), // LUT input
                .I1(in_1_i[87]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_86(.O(out[86]),     // LUT general output
                .I0(in_0_i[86]), // LUT input
                .I1(in_1_i[86]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_85(.O(out[85]),     // LUT general output
                .I0(in_0_i[85]), // LUT input
                .I1(in_1_i[85]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_84(.O(out[84]),     // LUT general output
                .I0(in_0_i[84]), // LUT input
                .I1(in_1_i[84]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_83(.O(out[83]),     // LUT general output
                .I0(in_0_i[83]), // LUT input
                .I1(in_1_i[83]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_82(.O(out[82]),     // LUT general output
                .I0(in_0_i[82]), // LUT input
                .I1(in_1_i[82]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_81(.O(out[81]),     // LUT general output
                .I0(in_0_i[81]), // LUT input
                .I1(in_1_i[81]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_80(.O(out[80]),     // LUT general output
                .I0(in_0_i[80]), // LUT input
                .I1(in_1_i[80]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_79(.O(out[79]),     // LUT general output
                .I0(in_0_i[79]), // LUT input
                .I1(in_1_i[79]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_78(.O(out[78]),     // LUT general output
                .I0(in_0_i[78]), // LUT input
                .I1(in_1_i[78]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_77(.O(out[77]),     // LUT general output
                .I0(in_0_i[77]), // LUT input
                .I1(in_1_i[77]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_76(.O(out[76]),     // LUT general output
                .I0(in_0_i[76]), // LUT input
                .I1(in_1_i[76]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_75(.O(out[75]),     // LUT general output
                .I0(in_0_i[75]), // LUT input
                .I1(in_1_i[75]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_74(.O(out[74]),     // LUT general output
                .I0(in_0_i[74]), // LUT input
                .I1(in_1_i[74]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_73(.O(out[73]),     // LUT general output
                .I0(in_0_i[73]), // LUT input
                .I1(in_1_i[73]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_72(.O(out[72]),     // LUT general output
                .I0(in_0_i[72]), // LUT input
                .I1(in_1_i[72]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_71(.O(out[71]),     // LUT general output
                .I0(in_0_i[71]), // LUT input
                .I1(in_1_i[71]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_70(.O(out[70]),     // LUT general output
                .I0(in_0_i[70]), // LUT input
                .I1(in_1_i[70]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_69(.O(out[69]),     // LUT general output
                .I0(in_0_i[69]), // LUT input
                .I1(in_1_i[69]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_68(.O(out[68]),     // LUT general output
                .I0(in_0_i[68]), // LUT input
                .I1(in_1_i[68]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_67(.O(out[67]),     // LUT general output
                .I0(in_0_i[67]), // LUT input
                .I1(in_1_i[67]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_66(.O(out[66]),     // LUT general output
                .I0(in_0_i[66]), // LUT input
                .I1(in_1_i[66]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_65(.O(out[65]),     // LUT general output
                .I0(in_0_i[65]), // LUT input
                .I1(in_1_i[65]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_64(.O(out[64]),     // LUT general output
                .I0(in_0_i[64]), // LUT input
                .I1(in_1_i[64]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_63(.O(out[63]),     // LUT general output
                .I0(in_0_i[63]), // LUT input
                .I1(in_1_i[63]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_62(.O(out[62]),     // LUT general output
                .I0(in_0_i[62]), // LUT input
                .I1(in_1_i[62]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_61(.O(out[61]),     // LUT general output
                .I0(in_0_i[61]), // LUT input
                .I1(in_1_i[61]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_60(.O(out[60]),     // LUT general output
                .I0(in_0_i[60]), // LUT input
                .I1(in_1_i[60]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_59(.O(out[59]),     // LUT general output
                .I0(in_0_i[59]), // LUT input
                .I1(in_1_i[59]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_58(.O(out[58]),     // LUT general output
                .I0(in_0_i[58]), // LUT input
                .I1(in_1_i[58]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_57(.O(out[57]),     // LUT general output
                .I0(in_0_i[57]), // LUT input
                .I1(in_1_i[57]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_56(.O(out[56]),     // LUT general output
                .I0(in_0_i[56]), // LUT input
                .I1(in_1_i[56]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_55(.O(out[55]),     // LUT general output
                .I0(in_0_i[55]), // LUT input
                .I1(in_1_i[55]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_54(.O(out[54]),     // LUT general output
                .I0(in_0_i[54]), // LUT input
                .I1(in_1_i[54]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_53(.O(out[53]),     // LUT general output
                .I0(in_0_i[53]), // LUT input
                .I1(in_1_i[53]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_52(.O(out[52]),     // LUT general output
                .I0(in_0_i[52]), // LUT input
                .I1(in_1_i[52]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_51(.O(out[51]),     // LUT general output
                .I0(in_0_i[51]), // LUT input
                .I1(in_1_i[51]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_50(.O(out[50]),     // LUT general output
                .I0(in_0_i[50]), // LUT input
                .I1(in_1_i[50]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_49(.O(out[49]),     // LUT general output
                .I0(in_0_i[49]), // LUT input
                .I1(in_1_i[49]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_48(.O(out[48]),     // LUT general output
                .I0(in_0_i[48]), // LUT input
                .I1(in_1_i[48]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_47(.O(out[47]),     // LUT general output
                .I0(in_0_i[47]), // LUT input
                .I1(in_1_i[47]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_46(.O(out[46]),     // LUT general output
                .I0(in_0_i[46]), // LUT input
                .I1(in_1_i[46]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_45(.O(out[45]),     // LUT general output
                .I0(in_0_i[45]), // LUT input
                .I1(in_1_i[45]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_44(.O(out[44]),     // LUT general output
                .I0(in_0_i[44]), // LUT input
                .I1(in_1_i[44]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_43(.O(out[43]),     // LUT general output
                .I0(in_0_i[43]), // LUT input
                .I1(in_1_i[43]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_42(.O(out[42]),     // LUT general output
                .I0(in_0_i[42]), // LUT input
                .I1(in_1_i[42]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_41(.O(out[41]),     // LUT general output
                .I0(in_0_i[41]), // LUT input
                .I1(in_1_i[41]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_40(.O(out[40]),     // LUT general output
                .I0(in_0_i[40]), // LUT input
                .I1(in_1_i[40]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_39(.O(out[39]),     // LUT general output
                .I0(in_0_i[39]), // LUT input
                .I1(in_1_i[39]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_38(.O(out[38]),     // LUT general output
                .I0(in_0_i[38]), // LUT input
                .I1(in_1_i[38]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_37(.O(out[37]),     // LUT general output
                .I0(in_0_i[37]), // LUT input
                .I1(in_1_i[37]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_36(.O(out[36]),     // LUT general output
                .I0(in_0_i[36]), // LUT input
                .I1(in_1_i[36]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_35(.O(out[35]),     // LUT general output
                .I0(in_0_i[35]), // LUT input
                .I1(in_1_i[35]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_34(.O(out[34]),     // LUT general output
                .I0(in_0_i[34]), // LUT input
                .I1(in_1_i[34]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_33(.O(out[33]),     // LUT general output
                .I0(in_0_i[33]), // LUT input
                .I1(in_1_i[33]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_32(.O(out[32]),     // LUT general output
                .I0(in_0_i[32]), // LUT input
                .I1(in_1_i[32]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_31(.O(out[31]),     // LUT general output
                .I0(in_0_i[31]), // LUT input
                .I1(in_1_i[31]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_30(.O(out[30]),     // LUT general output
                .I0(in_0_i[30]), // LUT input
                .I1(in_1_i[30]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_29(.O(out[29]),     // LUT general output
                .I0(in_0_i[29]), // LUT input
                .I1(in_1_i[29]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_28(.O(out[28]),     // LUT general output
                .I0(in_0_i[28]), // LUT input
                .I1(in_1_i[28]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_27(.O(out[27]),     // LUT general output
                .I0(in_0_i[27]), // LUT input
                .I1(in_1_i[27]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_26(.O(out[26]),     // LUT general output
                .I0(in_0_i[26]), // LUT input
                .I1(in_1_i[26]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_25(.O(out[25]),     // LUT general output
                .I0(in_0_i[25]), // LUT input
                .I1(in_1_i[25]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_24(.O(out[24]),     // LUT general output
                .I0(in_0_i[24]), // LUT input
                .I1(in_1_i[24]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_23(.O(out[23]),     // LUT general output
                .I0(in_0_i[23]), // LUT input
                .I1(in_1_i[23]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_22(.O(out[22]),     // LUT general output
                .I0(in_0_i[22]), // LUT input
                .I1(in_1_i[22]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_21(.O(out[21]),     // LUT general output
                .I0(in_0_i[21]), // LUT input
                .I1(in_1_i[21]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_20(.O(out[20]),     // LUT general output
                .I0(in_0_i[20]), // LUT input
                .I1(in_1_i[20]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_19(.O(out[19]),     // LUT general output
                .I0(in_0_i[19]), // LUT input
                .I1(in_1_i[19]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_18(.O(out[18]),     // LUT general output
                .I0(in_0_i[18]), // LUT input
                .I1(in_1_i[18]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_17(.O(out[17]),     // LUT general output
                .I0(in_0_i[17]), // LUT input
                .I1(in_1_i[17]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_16(.O(out[16]),     // LUT general output
                .I0(in_0_i[16]), // LUT input
                .I1(in_1_i[16]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_15(.O(out[15]),     // LUT general output
                .I0(in_0_i[15]), // LUT input
                .I1(in_1_i[15]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_14(.O(out[14]),     // LUT general output
                .I0(in_0_i[14]), // LUT input
                .I1(in_1_i[14]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_13(.O(out[13]),     // LUT general output
                .I0(in_0_i[13]), // LUT input
                .I1(in_1_i[13]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_12(.O(out[12]),     // LUT general output
                .I0(in_0_i[12]), // LUT input
                .I1(in_1_i[12]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_11(.O(out[11]),     // LUT general output
                .I0(in_0_i[11]), // LUT input
                .I1(in_1_i[11]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_10(.O(out[10]),     // LUT general output
                .I0(in_0_i[10]), // LUT input
                .I1(in_1_i[10]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_9(.O(out[9]),     // LUT general output
                .I0(in_0_i[9]), // LUT input
                .I1(in_1_i[9]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_8(.O(out[8]),     // LUT general output
                .I0(in_0_i[8]), // LUT input
                .I1(in_1_i[8]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_7(.O(out[7]),     // LUT general output
                .I0(in_0_i[7]), // LUT input
                .I1(in_1_i[7]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_6(.O(out[6]),     // LUT general output
                .I0(in_0_i[6]), // LUT input
                .I1(in_1_i[6]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_5(.O(out[5]),     // LUT general output
                .I0(in_0_i[5]), // LUT input
                .I1(in_1_i[5]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_4(.O(out[4]),     // LUT general output
                .I0(in_0_i[4]), // LUT input
                .I1(in_1_i[4]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_3(.O(out[3]),     // LUT general output
                .I0(in_0_i[3]), // LUT input
                .I1(in_1_i[3]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_2(.O(out[2]),     // LUT general output
                .I0(in_0_i[2]), // LUT input
                .I1(in_1_i[2]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_1(.O(out[1]),     // LUT general output
                .I0(in_0_i[1]), // LUT input
                .I1(in_1_i[1]), // LUT input
                .I2(sel_i)     // LUT input
          );
    LUT3 #(
                .INIT(8'hca)         // Specify LUT Contents
            )mux_0(.O(out[0]),     // LUT general output
                .I0(in_0_i[0]), // LUT input
                .I1(in_1_i[0]), // LUT input
                .I2(sel_i)     // LUT input
          );

endmodule
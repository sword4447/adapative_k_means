`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 05/12/2021 11:58:55 PM
// Design Name: 
// Module Name: mux_16i1o_32b_no_dly
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module mux_16i1o_32b_no_dly(
	input  [31:0]  din_0_i,
	input  [31:0]  din_1_i,
	input  [31:0]  din_2_i,
	input  [31:0]  din_3_i,	
	input  [31:0]  din_4_i,
	input  [31:0]  din_5_i,
	input  [31:0]  din_6_i,
	input  [31:0]  din_7_i,	 
	input  [31:0]  din_8_i,
	input  [31:0]  din_9_i,
	input  [31:0]  din_10_i,
	input  [31:0]  din_11_i,	
	input  [31:0]  din_12_i,
	input  [31:0]  din_13_i,
	input  [31:0]  din_14_i,
	input  [31:0]  din_15_i,	 	 

    input  [3:0]  sel_i,
	 
    output [31:0]  dout_o
    );
        Mux_16I1O_1b_no_dly dout_b31_inst (
    .din_0_i(din_0_i[31]),
     .din_1_i(din_1_i[31]),
     .din_2_i(din_2_i[31]),
    .din_3_i(din_3_i[31]),
    .din_4_i(din_4_i[31]),
     .din_5_i(din_5_i[31]),
    .din_6_i(din_6_i[31]),
     .din_7_i(din_7_i[31]),
    .din_8_i(din_8_i[31]),
    .din_9_i(din_9_i[31]),
     .din_10_i(din_10_i[31]),
    .din_11_i(din_11_i[31]),
     .din_12_i(din_12_i[31]),
    .din_13_i(din_13_i[31]),
    .din_14_i(din_14_i[31]),
    .din_15_i(din_15_i[31]),
    .sel_i(sel_i),
    .dout_o(dout_o[31])
    );
    Mux_16I1O_1b_no_dly dout_b30_inst (
    .din_0_i(din_0_i[30]),
     .din_1_i(din_1_i[30]),
     .din_2_i(din_2_i[30]),
    .din_3_i(din_3_i[30]),
    .din_4_i(din_4_i[30]),
     .din_5_i(din_5_i[30]),
    .din_6_i(din_6_i[30]),
     .din_7_i(din_7_i[30]),
    .din_8_i(din_8_i[30]),
    .din_9_i(din_9_i[30]),
     .din_10_i(din_10_i[30]),
    .din_11_i(din_11_i[30]),
     .din_12_i(din_12_i[30]),
    .din_13_i(din_13_i[30]),
    .din_14_i(din_14_i[30]),
    .din_15_i(din_15_i[30]),
    .sel_i(sel_i),
    .dout_o(dout_o[30])
    );
    Mux_16I1O_1b_no_dly dout_b29_inst (
    .din_0_i(din_0_i[29]),
     .din_1_i(din_1_i[29]),
     .din_2_i(din_2_i[29]),
    .din_3_i(din_3_i[29]),
    .din_4_i(din_4_i[29]),
     .din_5_i(din_5_i[29]),
    .din_6_i(din_6_i[29]),
     .din_7_i(din_7_i[29]),
    .din_8_i(din_8_i[29]),
    .din_9_i(din_9_i[29]),
     .din_10_i(din_10_i[29]),
    .din_11_i(din_11_i[29]),
     .din_12_i(din_12_i[29]),
    .din_13_i(din_13_i[29]),
    .din_14_i(din_14_i[29]),
    .din_15_i(din_15_i[29]),
    .sel_i(sel_i),
    .dout_o(dout_o[29])
    );
    Mux_16I1O_1b_no_dly dout_b28_inst (
    .din_0_i(din_0_i[28]),
     .din_1_i(din_1_i[28]),
     .din_2_i(din_2_i[28]),
    .din_3_i(din_3_i[28]),
    .din_4_i(din_4_i[28]),
     .din_5_i(din_5_i[28]),
    .din_6_i(din_6_i[28]),
     .din_7_i(din_7_i[28]),
    .din_8_i(din_8_i[28]),
    .din_9_i(din_9_i[28]),
     .din_10_i(din_10_i[28]),
    .din_11_i(din_11_i[28]),
     .din_12_i(din_12_i[28]),
    .din_13_i(din_13_i[28]),
    .din_14_i(din_14_i[28]),
    .din_15_i(din_15_i[28]),
    .sel_i(sel_i),
    .dout_o(dout_o[28])
    );
    Mux_16I1O_1b_no_dly dout_b27_inst (
    .din_0_i(din_0_i[27]),
     .din_1_i(din_1_i[27]),
     .din_2_i(din_2_i[27]),
    .din_3_i(din_3_i[27]),
    .din_4_i(din_4_i[27]),
     .din_5_i(din_5_i[27]),
    .din_6_i(din_6_i[27]),
     .din_7_i(din_7_i[27]),
    .din_8_i(din_8_i[27]),
    .din_9_i(din_9_i[27]),
     .din_10_i(din_10_i[27]),
    .din_11_i(din_11_i[27]),
     .din_12_i(din_12_i[27]),
    .din_13_i(din_13_i[27]),
    .din_14_i(din_14_i[27]),
    .din_15_i(din_15_i[27]),
    .sel_i(sel_i),
    .dout_o(dout_o[27])
    );
    Mux_16I1O_1b_no_dly dout_b26_inst (
    .din_0_i(din_0_i[26]),
     .din_1_i(din_1_i[26]),
     .din_2_i(din_2_i[26]),
    .din_3_i(din_3_i[26]),
    .din_4_i(din_4_i[26]),
     .din_5_i(din_5_i[26]),
    .din_6_i(din_6_i[26]),
     .din_7_i(din_7_i[26]),
    .din_8_i(din_8_i[26]),
    .din_9_i(din_9_i[26]),
     .din_10_i(din_10_i[26]),
    .din_11_i(din_11_i[26]),
     .din_12_i(din_12_i[26]),
    .din_13_i(din_13_i[26]),
    .din_14_i(din_14_i[26]),
    .din_15_i(din_15_i[26]),
    .sel_i(sel_i),
    .dout_o(dout_o[26])
    );
    Mux_16I1O_1b_no_dly dout_b25_inst (
    .din_0_i(din_0_i[25]),
     .din_1_i(din_1_i[25]),
     .din_2_i(din_2_i[25]),
    .din_3_i(din_3_i[25]),
    .din_4_i(din_4_i[25]),
     .din_5_i(din_5_i[25]),
    .din_6_i(din_6_i[25]),
     .din_7_i(din_7_i[25]),
    .din_8_i(din_8_i[25]),
    .din_9_i(din_9_i[25]),
     .din_10_i(din_10_i[25]),
    .din_11_i(din_11_i[25]),
     .din_12_i(din_12_i[25]),
    .din_13_i(din_13_i[25]),
    .din_14_i(din_14_i[25]),
    .din_15_i(din_15_i[25]),
    .sel_i(sel_i),
    .dout_o(dout_o[25])
    );
    Mux_16I1O_1b_no_dly dout_b24_inst (
    .din_0_i(din_0_i[24]),
     .din_1_i(din_1_i[24]),
     .din_2_i(din_2_i[24]),
    .din_3_i(din_3_i[24]),
    .din_4_i(din_4_i[24]),
     .din_5_i(din_5_i[24]),
    .din_6_i(din_6_i[24]),
     .din_7_i(din_7_i[24]),
    .din_8_i(din_8_i[24]),
    .din_9_i(din_9_i[24]),
     .din_10_i(din_10_i[24]),
    .din_11_i(din_11_i[24]),
     .din_12_i(din_12_i[24]),
    .din_13_i(din_13_i[24]),
    .din_14_i(din_14_i[24]),
    .din_15_i(din_15_i[24]),
    .sel_i(sel_i),
    .dout_o(dout_o[24])
    );
    Mux_16I1O_1b_no_dly dout_b23_inst (
    .din_0_i(din_0_i[23]),
     .din_1_i(din_1_i[23]),
     .din_2_i(din_2_i[23]),
    .din_3_i(din_3_i[23]),
    .din_4_i(din_4_i[23]),
     .din_5_i(din_5_i[23]),
    .din_6_i(din_6_i[23]),
     .din_7_i(din_7_i[23]),
    .din_8_i(din_8_i[23]),
    .din_9_i(din_9_i[23]),
     .din_10_i(din_10_i[23]),
    .din_11_i(din_11_i[23]),
     .din_12_i(din_12_i[23]),
    .din_13_i(din_13_i[23]),
    .din_14_i(din_14_i[23]),
    .din_15_i(din_15_i[23]),
    .sel_i(sel_i),
    .dout_o(dout_o[23])
    );
    Mux_16I1O_1b_no_dly dout_b22_inst (
    .din_0_i(din_0_i[22]),
     .din_1_i(din_1_i[22]),
     .din_2_i(din_2_i[22]),
    .din_3_i(din_3_i[22]),
    .din_4_i(din_4_i[22]),
     .din_5_i(din_5_i[22]),
    .din_6_i(din_6_i[22]),
     .din_7_i(din_7_i[22]),
    .din_8_i(din_8_i[22]),
    .din_9_i(din_9_i[22]),
     .din_10_i(din_10_i[22]),
    .din_11_i(din_11_i[22]),
     .din_12_i(din_12_i[22]),
    .din_13_i(din_13_i[22]),
    .din_14_i(din_14_i[22]),
    .din_15_i(din_15_i[22]),
    .sel_i(sel_i),
    .dout_o(dout_o[22])
    );
    Mux_16I1O_1b_no_dly dout_b21_inst (
    .din_0_i(din_0_i[21]),
     .din_1_i(din_1_i[21]),
     .din_2_i(din_2_i[21]),
    .din_3_i(din_3_i[21]),
    .din_4_i(din_4_i[21]),
     .din_5_i(din_5_i[21]),
    .din_6_i(din_6_i[21]),
     .din_7_i(din_7_i[21]),
    .din_8_i(din_8_i[21]),
    .din_9_i(din_9_i[21]),
     .din_10_i(din_10_i[21]),
    .din_11_i(din_11_i[21]),
     .din_12_i(din_12_i[21]),
    .din_13_i(din_13_i[21]),
    .din_14_i(din_14_i[21]),
    .din_15_i(din_15_i[21]),
    .sel_i(sel_i),
    .dout_o(dout_o[21])
    );
    Mux_16I1O_1b_no_dly dout_b20_inst (
    .din_0_i(din_0_i[20]),
     .din_1_i(din_1_i[20]),
     .din_2_i(din_2_i[20]),
    .din_3_i(din_3_i[20]),
    .din_4_i(din_4_i[20]),
     .din_5_i(din_5_i[20]),
    .din_6_i(din_6_i[20]),
     .din_7_i(din_7_i[20]),
    .din_8_i(din_8_i[20]),
    .din_9_i(din_9_i[20]),
     .din_10_i(din_10_i[20]),
    .din_11_i(din_11_i[20]),
     .din_12_i(din_12_i[20]),
    .din_13_i(din_13_i[20]),
    .din_14_i(din_14_i[20]),
    .din_15_i(din_15_i[20]),
    .sel_i(sel_i),
    .dout_o(dout_o[20])
    );
    Mux_16I1O_1b_no_dly dout_b19_inst (
    .din_0_i(din_0_i[19]),
     .din_1_i(din_1_i[19]),
     .din_2_i(din_2_i[19]),
    .din_3_i(din_3_i[19]),
    .din_4_i(din_4_i[19]),
     .din_5_i(din_5_i[19]),
    .din_6_i(din_6_i[19]),
     .din_7_i(din_7_i[19]),
    .din_8_i(din_8_i[19]),
    .din_9_i(din_9_i[19]),
     .din_10_i(din_10_i[19]),
    .din_11_i(din_11_i[19]),
     .din_12_i(din_12_i[19]),
    .din_13_i(din_13_i[19]),
    .din_14_i(din_14_i[19]),
    .din_15_i(din_15_i[19]),
    .sel_i(sel_i),
    .dout_o(dout_o[19])
    );
    Mux_16I1O_1b_no_dly dout_b18_inst (
    .din_0_i(din_0_i[18]),
     .din_1_i(din_1_i[18]),
     .din_2_i(din_2_i[18]),
    .din_3_i(din_3_i[18]),
    .din_4_i(din_4_i[18]),
     .din_5_i(din_5_i[18]),
    .din_6_i(din_6_i[18]),
     .din_7_i(din_7_i[18]),
    .din_8_i(din_8_i[18]),
    .din_9_i(din_9_i[18]),
     .din_10_i(din_10_i[18]),
    .din_11_i(din_11_i[18]),
     .din_12_i(din_12_i[18]),
    .din_13_i(din_13_i[18]),
    .din_14_i(din_14_i[18]),
    .din_15_i(din_15_i[18]),
    .sel_i(sel_i),
    .dout_o(dout_o[18])
    );
    Mux_16I1O_1b_no_dly dout_b17_inst (
    .din_0_i(din_0_i[17]),
     .din_1_i(din_1_i[17]),
     .din_2_i(din_2_i[17]),
    .din_3_i(din_3_i[17]),
    .din_4_i(din_4_i[17]),
     .din_5_i(din_5_i[17]),
    .din_6_i(din_6_i[17]),
     .din_7_i(din_7_i[17]),
    .din_8_i(din_8_i[17]),
    .din_9_i(din_9_i[17]),
     .din_10_i(din_10_i[17]),
    .din_11_i(din_11_i[17]),
     .din_12_i(din_12_i[17]),
    .din_13_i(din_13_i[17]),
    .din_14_i(din_14_i[17]),
    .din_15_i(din_15_i[17]),
    .sel_i(sel_i),
    .dout_o(dout_o[17])
    );
    Mux_16I1O_1b_no_dly dout_b16_inst (
    .din_0_i(din_0_i[16]),
     .din_1_i(din_1_i[16]),
     .din_2_i(din_2_i[16]),
    .din_3_i(din_3_i[16]),
    .din_4_i(din_4_i[16]),
     .din_5_i(din_5_i[16]),
    .din_6_i(din_6_i[16]),
     .din_7_i(din_7_i[16]),
    .din_8_i(din_8_i[16]),
    .din_9_i(din_9_i[16]),
     .din_10_i(din_10_i[16]),
    .din_11_i(din_11_i[16]),
     .din_12_i(din_12_i[16]),
    .din_13_i(din_13_i[16]),
    .din_14_i(din_14_i[16]),
    .din_15_i(din_15_i[16]),
    .sel_i(sel_i),
    .dout_o(dout_o[16])
    );
    Mux_16I1O_1b_no_dly dout_b15_inst (
    .din_0_i(din_0_i[15]),
     .din_1_i(din_1_i[15]),
     .din_2_i(din_2_i[15]),
    .din_3_i(din_3_i[15]),
    .din_4_i(din_4_i[15]),
     .din_5_i(din_5_i[15]),
    .din_6_i(din_6_i[15]),
     .din_7_i(din_7_i[15]),
    .din_8_i(din_8_i[15]),
    .din_9_i(din_9_i[15]),
     .din_10_i(din_10_i[15]),
    .din_11_i(din_11_i[15]),
     .din_12_i(din_12_i[15]),
    .din_13_i(din_13_i[15]),
    .din_14_i(din_14_i[15]),
    .din_15_i(din_15_i[15]),
    .sel_i(sel_i),
    .dout_o(dout_o[15])
    );
    Mux_16I1O_1b_no_dly dout_b14_inst (
    .din_0_i(din_0_i[14]),
     .din_1_i(din_1_i[14]),
     .din_2_i(din_2_i[14]),
    .din_3_i(din_3_i[14]),
    .din_4_i(din_4_i[14]),
     .din_5_i(din_5_i[14]),
    .din_6_i(din_6_i[14]),
     .din_7_i(din_7_i[14]),
    .din_8_i(din_8_i[14]),
    .din_9_i(din_9_i[14]),
     .din_10_i(din_10_i[14]),
    .din_11_i(din_11_i[14]),
     .din_12_i(din_12_i[14]),
    .din_13_i(din_13_i[14]),
    .din_14_i(din_14_i[14]),
    .din_15_i(din_15_i[14]),
    .sel_i(sel_i),
    .dout_o(dout_o[14])
    );
    Mux_16I1O_1b_no_dly dout_b13_inst (
    .din_0_i(din_0_i[13]),
     .din_1_i(din_1_i[13]),
     .din_2_i(din_2_i[13]),
    .din_3_i(din_3_i[13]),
    .din_4_i(din_4_i[13]),
     .din_5_i(din_5_i[13]),
    .din_6_i(din_6_i[13]),
     .din_7_i(din_7_i[13]),
    .din_8_i(din_8_i[13]),
    .din_9_i(din_9_i[13]),
     .din_10_i(din_10_i[13]),
    .din_11_i(din_11_i[13]),
     .din_12_i(din_12_i[13]),
    .din_13_i(din_13_i[13]),
    .din_14_i(din_14_i[13]),
    .din_15_i(din_15_i[13]),
    .sel_i(sel_i),
    .dout_o(dout_o[13])
    );
    Mux_16I1O_1b_no_dly dout_b12_inst (
    .din_0_i(din_0_i[12]),
     .din_1_i(din_1_i[12]),
     .din_2_i(din_2_i[12]),
    .din_3_i(din_3_i[12]),
    .din_4_i(din_4_i[12]),
     .din_5_i(din_5_i[12]),
    .din_6_i(din_6_i[12]),
     .din_7_i(din_7_i[12]),
    .din_8_i(din_8_i[12]),
    .din_9_i(din_9_i[12]),
     .din_10_i(din_10_i[12]),
    .din_11_i(din_11_i[12]),
     .din_12_i(din_12_i[12]),
    .din_13_i(din_13_i[12]),
    .din_14_i(din_14_i[12]),
    .din_15_i(din_15_i[12]),
    .sel_i(sel_i),
    .dout_o(dout_o[12])
    );
    Mux_16I1O_1b_no_dly dout_b11_inst (
    .din_0_i(din_0_i[11]),
     .din_1_i(din_1_i[11]),
     .din_2_i(din_2_i[11]),
    .din_3_i(din_3_i[11]),
    .din_4_i(din_4_i[11]),
     .din_5_i(din_5_i[11]),
    .din_6_i(din_6_i[11]),
     .din_7_i(din_7_i[11]),
    .din_8_i(din_8_i[11]),
    .din_9_i(din_9_i[11]),
     .din_10_i(din_10_i[11]),
    .din_11_i(din_11_i[11]),
     .din_12_i(din_12_i[11]),
    .din_13_i(din_13_i[11]),
    .din_14_i(din_14_i[11]),
    .din_15_i(din_15_i[11]),
    .sel_i(sel_i),
    .dout_o(dout_o[11])
    );
    Mux_16I1O_1b_no_dly dout_b10_inst (
    .din_0_i(din_0_i[10]),
     .din_1_i(din_1_i[10]),
     .din_2_i(din_2_i[10]),
    .din_3_i(din_3_i[10]),
    .din_4_i(din_4_i[10]),
     .din_5_i(din_5_i[10]),
    .din_6_i(din_6_i[10]),
     .din_7_i(din_7_i[10]),
    .din_8_i(din_8_i[10]),
    .din_9_i(din_9_i[10]),
     .din_10_i(din_10_i[10]),
    .din_11_i(din_11_i[10]),
     .din_12_i(din_12_i[10]),
    .din_13_i(din_13_i[10]),
    .din_14_i(din_14_i[10]),
    .din_15_i(din_15_i[10]),
    .sel_i(sel_i),
    .dout_o(dout_o[10])
    );
    Mux_16I1O_1b_no_dly dout_b9_inst (
    .din_0_i(din_0_i[9]),
     .din_1_i(din_1_i[9]),
     .din_2_i(din_2_i[9]),
    .din_3_i(din_3_i[9]),
    .din_4_i(din_4_i[9]),
     .din_5_i(din_5_i[9]),
    .din_6_i(din_6_i[9]),
     .din_7_i(din_7_i[9]),
    .din_8_i(din_8_i[9]),
    .din_9_i(din_9_i[9]),
     .din_10_i(din_10_i[9]),
    .din_11_i(din_11_i[9]),
     .din_12_i(din_12_i[9]),
    .din_13_i(din_13_i[9]),
    .din_14_i(din_14_i[9]),
    .din_15_i(din_15_i[9]),
    .sel_i(sel_i),
    .dout_o(dout_o[9])
    );
    Mux_16I1O_1b_no_dly dout_b8_inst (
    .din_0_i(din_0_i[8]),
     .din_1_i(din_1_i[8]),
     .din_2_i(din_2_i[8]),
    .din_3_i(din_3_i[8]),
    .din_4_i(din_4_i[8]),
     .din_5_i(din_5_i[8]),
    .din_6_i(din_6_i[8]),
     .din_7_i(din_7_i[8]),
    .din_8_i(din_8_i[8]),
    .din_9_i(din_9_i[8]),
     .din_10_i(din_10_i[8]),
    .din_11_i(din_11_i[8]),
     .din_12_i(din_12_i[8]),
    .din_13_i(din_13_i[8]),
    .din_14_i(din_14_i[8]),
    .din_15_i(din_15_i[8]),
    .sel_i(sel_i),
    .dout_o(dout_o[8])
    );
    Mux_16I1O_1b_no_dly dout_b7_inst (
    .din_0_i(din_0_i[7]),
     .din_1_i(din_1_i[7]),
     .din_2_i(din_2_i[7]),
    .din_3_i(din_3_i[7]),
    .din_4_i(din_4_i[7]),
     .din_5_i(din_5_i[7]),
    .din_6_i(din_6_i[7]),
     .din_7_i(din_7_i[7]),
    .din_8_i(din_8_i[7]),
    .din_9_i(din_9_i[7]),
     .din_10_i(din_10_i[7]),
    .din_11_i(din_11_i[7]),
     .din_12_i(din_12_i[7]),
    .din_13_i(din_13_i[7]),
    .din_14_i(din_14_i[7]),
    .din_15_i(din_15_i[7]),
    .sel_i(sel_i),
    .dout_o(dout_o[7])
    );
    Mux_16I1O_1b_no_dly dout_b6_inst (
    .din_0_i(din_0_i[6]),
     .din_1_i(din_1_i[6]),
     .din_2_i(din_2_i[6]),
    .din_3_i(din_3_i[6]),
    .din_4_i(din_4_i[6]),
     .din_5_i(din_5_i[6]),
    .din_6_i(din_6_i[6]),
     .din_7_i(din_7_i[6]),
    .din_8_i(din_8_i[6]),
    .din_9_i(din_9_i[6]),
     .din_10_i(din_10_i[6]),
    .din_11_i(din_11_i[6]),
     .din_12_i(din_12_i[6]),
    .din_13_i(din_13_i[6]),
    .din_14_i(din_14_i[6]),
    .din_15_i(din_15_i[6]),
    .sel_i(sel_i),
    .dout_o(dout_o[6])
    );
    Mux_16I1O_1b_no_dly dout_b5_inst (
    .din_0_i(din_0_i[5]),
     .din_1_i(din_1_i[5]),
     .din_2_i(din_2_i[5]),
    .din_3_i(din_3_i[5]),
    .din_4_i(din_4_i[5]),
     .din_5_i(din_5_i[5]),
    .din_6_i(din_6_i[5]),
     .din_7_i(din_7_i[5]),
    .din_8_i(din_8_i[5]),
    .din_9_i(din_9_i[5]),
     .din_10_i(din_10_i[5]),
    .din_11_i(din_11_i[5]),
     .din_12_i(din_12_i[5]),
    .din_13_i(din_13_i[5]),
    .din_14_i(din_14_i[5]),
    .din_15_i(din_15_i[5]),
    .sel_i(sel_i),
    .dout_o(dout_o[5])
    );
    Mux_16I1O_1b_no_dly dout_b4_inst (
    .din_0_i(din_0_i[4]),
     .din_1_i(din_1_i[4]),
     .din_2_i(din_2_i[4]),
    .din_3_i(din_3_i[4]),
    .din_4_i(din_4_i[4]),
     .din_5_i(din_5_i[4]),
    .din_6_i(din_6_i[4]),
     .din_7_i(din_7_i[4]),
    .din_8_i(din_8_i[4]),
    .din_9_i(din_9_i[4]),
     .din_10_i(din_10_i[4]),
    .din_11_i(din_11_i[4]),
     .din_12_i(din_12_i[4]),
    .din_13_i(din_13_i[4]),
    .din_14_i(din_14_i[4]),
    .din_15_i(din_15_i[4]),
    .sel_i(sel_i),
    .dout_o(dout_o[4])
    );
    Mux_16I1O_1b_no_dly dout_b3_inst (
    .din_0_i(din_0_i[3]),
     .din_1_i(din_1_i[3]),
     .din_2_i(din_2_i[3]),
    .din_3_i(din_3_i[3]),
    .din_4_i(din_4_i[3]),
     .din_5_i(din_5_i[3]),
    .din_6_i(din_6_i[3]),
     .din_7_i(din_7_i[3]),
    .din_8_i(din_8_i[3]),
    .din_9_i(din_9_i[3]),
     .din_10_i(din_10_i[3]),
    .din_11_i(din_11_i[3]),
     .din_12_i(din_12_i[3]),
    .din_13_i(din_13_i[3]),
    .din_14_i(din_14_i[3]),
    .din_15_i(din_15_i[3]),
    .sel_i(sel_i),
    .dout_o(dout_o[3])
    );
    Mux_16I1O_1b_no_dly dout_b2_inst (
    .din_0_i(din_0_i[2]),
     .din_1_i(din_1_i[2]),
     .din_2_i(din_2_i[2]),
    .din_3_i(din_3_i[2]),
    .din_4_i(din_4_i[2]),
     .din_5_i(din_5_i[2]),
    .din_6_i(din_6_i[2]),
     .din_7_i(din_7_i[2]),
    .din_8_i(din_8_i[2]),
    .din_9_i(din_9_i[2]),
     .din_10_i(din_10_i[2]),
    .din_11_i(din_11_i[2]),
     .din_12_i(din_12_i[2]),
    .din_13_i(din_13_i[2]),
    .din_14_i(din_14_i[2]),
    .din_15_i(din_15_i[2]),
    .sel_i(sel_i),
    .dout_o(dout_o[2])
    );
    Mux_16I1O_1b_no_dly dout_b1_inst (
    .din_0_i(din_0_i[1]),
     .din_1_i(din_1_i[1]),
     .din_2_i(din_2_i[1]),
    .din_3_i(din_3_i[1]),
    .din_4_i(din_4_i[1]),
     .din_5_i(din_5_i[1]),
    .din_6_i(din_6_i[1]),
     .din_7_i(din_7_i[1]),
    .din_8_i(din_8_i[1]),
    .din_9_i(din_9_i[1]),
     .din_10_i(din_10_i[1]),
    .din_11_i(din_11_i[1]),
     .din_12_i(din_12_i[1]),
    .din_13_i(din_13_i[1]),
    .din_14_i(din_14_i[1]),
    .din_15_i(din_15_i[1]),
    .sel_i(sel_i),
    .dout_o(dout_o[1])
    );
    Mux_16I1O_1b_no_dly dout_b0_inst (
    .din_0_i(din_0_i[0]),
     .din_1_i(din_1_i[0]),
     .din_2_i(din_2_i[0]),
    .din_3_i(din_3_i[0]),
    .din_4_i(din_4_i[0]),
     .din_5_i(din_5_i[0]),
    .din_6_i(din_6_i[0]),
     .din_7_i(din_7_i[0]),
    .din_8_i(din_8_i[0]),
    .din_9_i(din_9_i[0]),
     .din_10_i(din_10_i[0]),
    .din_11_i(din_11_i[0]),
     .din_12_i(din_12_i[0]),
    .din_13_i(din_13_i[0]),
    .din_14_i(din_14_i[0]),
    .din_15_i(din_15_i[0]),
    .sel_i(sel_i),
    .dout_o(dout_o[0])
    );
endmodule
